��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a�����/�	v�+����@ɧ-3�����Iz�t�܀Le'H>	6"�U{��9�bEɤ6-�!�V��s� ���m�|����~μn���}�iԹ*VC�4���m7���-� �7�o�d�0w1 �⹺�)=k�:+5:� _M�e�$�"��O��0U̅�iZ��x�K�~̏*���;��R+X�="+$Y~�ml���n�H���K1,���0�ϔ���憲e'oN��D_lxY��^PZ�#�C�e��Au�֝��2ɤZ2���ܵ� �o���ǣߜM0ځr5r`D.ɩ�
e���
�Dc�����gC�8$����lc'�'@��A��Se��J�oY�\�?f�ᕭ�o0�\�O��H�$���m���M2�M��J��?�c��ˈA���~=ɮ�����D���B�p��;�e㹽yU4-����_8����p�R�C7�H��;v��F��5	��zMV�I�xB�cȀ�j��� l�{�I�e>;�IT�NF.v2���hb�]%fzy�0���#�%�GNאsXU�թ���*��j�5x
�P2V�?��9}��=�->���x�/#v��_�����J�N�(��x�USy��i7�4��J�ÞQb���u����V��i/��R�	J�,W��r����tx�E�r}ӣ��בrl��P=��������1+�&r�W]�#'`��5]h�?�G�i��:b�P�Ǎ�;�׈6����r�R�����
m;��V�j�w��^Q�Z1�d�p#��`�h� ����Ҹ"���'�1��o�}��d_��0�^$-9S������b�I'Ѿ(==� �����N^X39޻f�z�M߶�>m�84�G�d�|6� >��2'[�a[g� �oL�(Y�h/G���ܚ�ղy)a���l��� �d�,�f5�gFS4|�M8l> �����0<O`q�`�U�X�$.?@�S�xm���h*#���_��)��a��i��<g��Mە�����3xt�F�����ef̌�����:Pn�� EM�é�=����/�̣S1��$��<a��\u�!/�\����փ ���:�u���־��Q��2�sƴF�X�������)|=ZϠI�2É3�K�%3ń��q�؍o* t"it`�+��7��܌�G\{�ףm�8�~��#���hT���S-���@r��{�{�p�/��1�ȅ�M�J,��I�H��t��t+���z�ܤA�*?�����bW.���Jށh� 7J��5��T����ֽr�E7�����@n�KS+ư�pnT��s.��q0撍8f.x
�4��P��;��i�3�ԣ�@�}��)Z2��86��!R��.QL@`uJ%��л���"�T�o���4��t������������8]��T���]X{�;-|{�3���я�9&�D�ƞ~mt��L��d>��G}��P}�92��6�mhm��3�%������ڮ�e�v#V%|�Y�-F��I$S$���0��({O#SĂ��)'P>�Z"?�:H����2nȯvk�=�m�K�RT=9���IFsnVd	&��N!O.�3�o��-�5�����H�kc!tr��h�-��Ì����m��װ>g���i<ى�"�eNT�ؚ3�-q���H��ꦼ�����F�q�b��2f*�G)��>G�n�O��T�Lb&�,y� �w[�0�euDym��"�$�*����,�.�G�]��?��`�G\ɧ�N��>���t����T�K�E��cLM�^���%Tb��k���Bjth�++���}\f����[;vP<f��/[��B���f��>a�Ű���Pl��pް�.�_΄��e��,�ܮ5�=rT�/oܭ�Y� ��w���Kԅ�p$�h �A��Q|��d21��*���ѷmu���Jy��4u=3��۵T�@��(p���k�_�9�e�k �_��5��fK��
=�#h�g)��u�Z�b\��y���3��\=Hz�3�4D���"�!b��j�O������n(�%��eJ}Y`�}���خ����]݁���x�� w�)�0e�{���'B��l�m-�qkbM��ŵϭl��n-�C˼��,�ۓ�N�ń��ͬb�E�wX��ԆȄCP�Q]�]�P�^֫��:��A�����q` ������ob�כҦ��ygPo�d�A�5��)^�Y��"z�q��e�?���4)�W����W�V䇚�%��Q�r�
,�yr?�r�lt�q���ے�n�jg�Պ����?�^�rq�7l҆$\��?
��>���1Zb>.1���!C�����8��%�8:E��F�0�&b#=��\�d҃�NS;��;GN!(|k�h� :����BB�l@>_K˸Ru7#��(����{���_5���VF���dU�':5��o*�V,_�ah Sc7�&��nvqm�n���jq#7��|W�0Eñk�n�`�'���_ �Q�l���� Փs�g��K+Y� 7Zo����(��ض��Qj�!�2���3��\?��)��C��M[���9Z�Ί�dȾ�U`�oyյ�`�~�[�iΦd�A�C�(Ea2��z�1�L��P�v�s���A���׬^m`���o�������6�qخ��3�D��
�P�&������>����y|�ѝ'���C��o�qC��H��er�!�1{К)lFc3X��D���u:�Yc'��ҽ��B���g�Nl�f@��q�h��A���ޝ�:�CP��}|�m�0Y�Z6�nʏe�0r��u�Zf�޸I�cy�MFҩc�iv�P1�G|�
w�I��K�rz�%d���D�٤c�v54R�Q�� ����p'y%^��)]j.q^��t�����QË�"l������I�j���'?���P����hGRQ�	�����=�To��f7�����ѣ\���ꄭ���%CJw�\�-��0HJ>��m%����5'���^`ese����8�y�َ�h��t��|s���(�_����"�'�Z������P��	l�.��s�8��:��e��Z�8~��'ʵ/�2�/���n~�ׂS��8�2�r��:���Pq�2袜u�|{ȼ�.�A�����;+�Kz�.����ⲻE����@oqr�1{�N|B]i{n�^��,�Sb��1�����DmƤ���T�m��L��I�V��gP��,�����$���7@����qە�h�9ҕ^0U�#|�<��
�16f��6a���=eQ�����&?Pq�����k3�KՂ�c�^�x�6�`����!I����[�d �f�7��;����������-��E���d���@�F��tW=�������_�:?���'E�%y��c���$�ƒ�s̗+{��JS����_۰��$yC��(���#��>%r����F��� ��<?�n�$x6=߾�
�
K%�����0Ɏq݅x��]|I5���u:y�; �QH8D��M�&3uJ����_#3�K�N��͢	s�eb�V:���Ǆ`}�a�^�iբZ��C�M"�P7�qT�	�N�.��O�Z�U�b���)R�2	i'�%L�N�D�Q�4<�y^�i~�7�)��*O�k� �؄�����V.X�.��'@�����#\���79�~ο%_�Dn�;H����ۚՐ&����ֈr�H8)��:1��XPڇPC����R�t�z�h��Qޭ�Ъ�I-kxv9�P%ue+��%�2д�a�ZU�e���dW���@9�hV�tȵ��^E�j�'��$�/�DW{/��+�fS$�!�Qx]0`��4�eT?�s���ø("�*/�湞�	?�L����M]�w�9'����]:ac	�G���������]��p[o���;�tti�h�.P�T�`=1���pˍ�nm1T
	����'�z��d��(A���2~ ib$j�zl6+�����7D���K~1��ץ�D�߂�c�x��Xn��k�]����l��9U�T�jy�i��o����iaDZ�g-\wѾVC<�R�X�� (ր �	�e���%ȥ�À=����6�R�"pj���YyAn�0�c�#꼑���2�;]z�Vx�1N*ˍ��)�w��B���gL=��p�`1�m���~�DL9!W���h���L/�)�r_���8D�-��e�O�{�^��E!�g�v�v�]��>?t�5A7+���������Q�/��Ȳ�h��>6 ��H��]seq���0_9�l��ɦ��bk�;�LȘ��'�
�S�0�ȼJ8�MX���2O�>���&21�e�Y��_�<]0�Ɗ�T��`P����6\��(&8�+�ySlr-�<�r����s���p� ���z�t��"+�Ԕ�i���,i"UQp}�<�+�(��vp'bu�K�SI��J�UQ�Y��l�6XL��u���๐�X���_��%�$����	���@��~��sp� �E�����>��1K��ۛ�q�����n.d��ڴ`�3#���!����4s.�h'機��DM�V��.���F��Q�q����%�@�֒���|u�,�n�U� �������t���%/J��_p'*?��K"�exAW}��ciy���|w�4a��Y-�(�ENe��Z[8�BKTl�{(��o $^�f��!�r2�A7~��޼�R;u���L{`
�t(<�.(�T�;1��������s�;1�r���K�[0=l@v��u��� ���6Q^ۇB��G� �V�/0I��mNj��3CZ�yg�ms���vD�.0���H��@G�����M~r8j�����#���è�	�S�^h��Ȩ�]��Q8qE��.��k�}A��(�8�l $��7��K �zَ�ݬ1��C����σ�$ #��7̓�/}�m�*FUc�O���ߴ�Qؿ%yy[.�2�u,<�I䘄!�A�q�_�I��[؃�.���|"zE���������f<��q��e*����ę+�{9�_��H�-��&F�?����%l���k��R�y�4HC<Kh�3��9����<�X$w^�(?����G�>|U"}x���o���hѱ@��#5D��>��V��
��*�Mxl/��������'!�<�����y����iη�
���m˶��lE^onM0�}�Pn�^��^��*hE�Q��t�[�^��Gهy��Sc��_�բ�d��1Խ��,��g�=*	bp;s��)�vp�yF�v����mT��Gj�Q�F� ���A�_&w���fᘂ����/Ѩ��Q�$��4%W&HL�8;z�-ظ�+Y~o�o�A%����z���
�@����O\��i��#�����]��J��kw�r��	�y�ʹ̉F����3�����}���j������]f����IF���|ʍ��c�vX�"V7��3�c�màH�^���+9ʅ�pT�&�Hޢk�@
��o�+�"{̳�Vf@ʼ�i�|�[�9�w(06=9���X �a]{#�S�B���"���Ǔ�ڠ�*��zi��6�9��Փ��I!�Q�}4Djw�GZ*>�Y9�,�]eY�ѯ8Rc�FBl�g���o����.j�14(Z|e޾�^�<�k	F�I���of��p��/��7FZ��t������(M��׋gc���(x�X���ֽ_A;�ZՓ��8�
(�d�����獃���i%��;ԧ%סH��s{�D;㕠F�l#�9��!�8	�A>�u o�o��w���F�a��#Dd��vDi@{�A�P&��lʃ�F�PTeF5T����O�՘-���E�0�F#�S��R��Ϫ朵e�������@e�~�0d�7Z��MW���ou��<X6�:�m��t��@0��f��P�N��h��������_��2�9�A��to[Z¬�?���iDW�J0C?���_l.��L��Q� 2�ݏvnO:"��K��n�2+����nꢁ��"X���Ag9�A����{F��(�;0~k���蛈1f(���|�{�'M2���T��Z�(+�n�}����K�x���.h��|;�2$"�e��=���ý��Eâ5�yޯ�����r�7-Ŗ"Iv��[�۠v�m<��h�8Z�v*��=j��ܣ��&���=�B������Z�4�	��OM�'( ���cG$ʁ��u�p�[ ޖ �5�F�t0����E���f���R��8�mv<Q #�>�>hƛh�V�ҭ��J�`��%7�Aŀ:�0�<uM1��&'�$	�Їy��40u�P�����	zHߣ�{%xJQy�ē��s��� �[�N��U���ΰIc�ϥl�������g'�S� "-���Ό-a�'ѝv�d8na��: �3�ǎ+ �鶴n���A�r!ܗ�"�fӪ�$$jQ�Ο��d���y9XsD�����,��3�p�/�"5y��66�+Y*�E������C�S�BcC٠_B��Տԙ���V���ậ�/_'y%y�uG��;����!�Rc���ޝ8�����d �t��A\F1xuub%����p;j��nX�!�~��w����/य़ ��b��������Խ�v"�(:�!T�q\'��}������s����� ��0]�\G��eV}z�	�`�D�Z�'�^���iP���Ε��a��D�awi��ǧ�n�&u�)�I~��;����%
��^*F�h"��-��j��j �������y&��ˈO�(B�U�ɓ���n�$3�vf�+m�+,0�h�P9�ӣ}Y7!�^�sD6���}�v����BI%��P�0�
2�s
��T��@���OS���7��֚�
+gA��	^u�=4Ȧ��%��w��Fp�N<�>2:ї�W5����l�x2�iA����4�D@����0�����_�"���������@CdQNe2j6ｊ�۝y'Vͺ�Hi���rs�'��
l2��;��Aze�D�#/����6��mזRK1.�Z�S4��$A%:΅�b������u��=��[N(����:�Y��Z����E������i�Ew��Y���'2_fH���S��s�~�#:8��AbI��E�+e�&����A{Ѿ������%�H��n]��
O��*~L�x,�_'���#yA�:'�k>����i�#��j��b�opD�+�]�h?��~4ˏo<Z|y+�7�t���뽘"p3�
t��Q���Z������
�T	�-�%�9��u��+V���/��UG�01CF��3V����j���<o��@r|�Δ�-�������lǭz��d~	 �f�c�Q��R�;�;~or�/�=�P�G����n�AJ	&Ǒ�:����뎷I8��I?EE�6�7�7�� 4wM��iS��k�g��@����>�`Og�|o�9�N�2B��܍�Q5(8xN!�mͷخz�9�s�7��Gia��y�J�z7��X]��+���Y�ZD��hHE�IY7W}5�Qш3SpHS�Ԃ�e�<X%�n.���"$6џo�k� �Wkv���
�DPg����dR���]�-+���>��b�e������e��'N�(=b��!G2�'oB)K�O@�#a: K�ދf����s������\��t�1�RЗS1mQFR����:	*��#o�VT�bw����<d��*o��k�b�EA�Nn�e�����KZX�!��:*�p���d�&�oc:>m`6���9�k����Գ�2/�?Iy��ت�Kj8�9X׆�<A�e��TĤ�8w3�O���k@�49p��!cEJ޾O����\�/����]��CX��X>h�N�jHKߓ��{����3��,'XYA��Ӝ�f_������K9�Ի�����)ܡ����	1|�r[|!��F9N�W���J�gCpj �r������57A���>:��`�_�l�w�'3�=�� ����}�|Ie�%^�h��4�0O]�XZ@�I�e�|���Ŧ׷�]��
��t4�������h`�����BX�N4]i|��u���l�.{ӕ_�N��͏�!AJ^�|�+&���p��t�"�����B���D��%|,�%��� ̴�UHVy RyF_OCA�PS:P�ID�9�u��5�%��<;�N�(N�	�����a��7�aT$u����2�S�l�dW m��V��"�𨣩�>*,V� U�?΁� ��3r8�{{�e�\����Y������/�n�C�TU��2�ƶ��LG����q�_hڬ$U/�'��k�����|~0q�Ʈ�O)`R/�Ͻycu�M�J�nWͱ��/\�͕�KF�����N��;���B�G��{�aêU�����īx[.Ҥ9:PUk��v�jҲT��it����,zb�g/C
�~�L0+�펌zBv�JqF/Q��{��I�4���D�Y�񯩱�MI6*k'Ò���!��S�"a�&��ym���s)E� c�ҵ�y��s��~��p��-e��wL.`���������+�d<����c+����H`�'�՘.�qѥX�xUkX��b�#}�����"������	�	��
��U�e@%��e��MK����"�9��������)�����H��@HA��XIEnj�`E��7%�������:&����G_;� 5:�q��Yz �5�<�
(㸓a�m����'ya~\b��Ȃ�ppyB�
�-ב��������a���0d���³��INV��$�Er۫����k����\C"�@X"oJڦR����/���"� � eB�y-��dS�\�wx�@���?U�Ft�ݧ�� �TN�д:>Q{�8q�b��}��i������6*�gcu�lX]o连��FV喿��ʏ��2W�R���x�Մ��Q��������ZŶ6Z�s�x1��P�d��ÄQ�<&?�.؋F�E����HE��a҂�R羡7^U1��	�m���Heβ��lu�p����/K �XΙ�
y��SU��[��n���_���hj9p���0X$v�G�Bd�aXٖ6�}���6�XsY~�s��\�q���ky�%���D�@N�E}Ԯ���a�k x_�8�i�+��	=�$��XJ�K�����a*�����!FՑ�k�1���+HvnQ�xH"�8�Օ��۹�����K�.^z��2���^��;REu���^�O�g�l͛�Ŗ��X��X_����#a`x����g��@gr%a~�llj-0���*��ES\h�1T����Fx�yy�FjM���x�������.ʮ�c�o"�ɡ�f������V�[�r%j�ߙ�#ڶ�N�dO�H���ǹ�fo�k�	Jђ�����WQ���^s�}T�"���mXc���Pl��XV�̵�ܕS��<�&?��<M��i����#:J���#��6��I�>��ܛEbz�rn�W6p�aRd�ZNI������h%�0��ʥ��ēx�[�\����YI�9�s���;s�z<;����;/Y����>�+�EB���
��,�� cZ�{i0w³�4�Ƙ�yA�h[��Z�>����� �ȧ)��HY��xZ�h\D$�C%���P�+��ڗ%<�	�J�/@�%�q]\����3ńǙ��"�<��E������v�-�&��ݸ%�X,�gTh2�ғd�(m��G;߬���؄an�n�c(�gg��nc�����p�r��:�k�*MW��jm"��u�����EGQ��@�T�^g���j�l���Wl �T�Y@���]Z�f��� |t��s���?�x���>E���ܦlXh��K9>?��sڒ��]h[�g�Y�о��'��ƀ���`z+��P���|k�2�ؕV18�Ƽ0IPB[˗��N��?� �� �b%@�q�/�G��,2M�*�f�/������O1��,��	L�֜'�~��ͻĤ i�^|Oqŗſ�w�W�Ƞ(���������J|����¢s��2�ʖf-j�������P��@��o"��4g�(Z=)�?$ۗ~9A�~!H2=C�ͅ�k�p9�p��+�I]�R���k�7��1�P)$�;�u[�P�kCS@R/&J?�͐�ih�mUBjy�=Y&�jDТ�޽��0<����6ƶ�y��D��AtD8ț�ԧ�5Shl
���ff���F����� � ���3	~�J2J�&�=N���.�8� �$Q�S��a/�}��3�P��Vh\�6�o ��2�t��y�o���b����1޷6�b��q3��f{�����϶6�ؚ�:�����̟��v�|�f�~f��|p�lI/��u�%7u��=��m��?�:F[��"@�����v���z��#�R������'���B���D�|�L�ё�ėj�Ac��B|G��c���1�t���]|��D���8���ѿ]yV|���
��~��k�ozś!���ko�*�r�g綄�&DX�1@��w<��L�a><xPp�T�N4z����'FR-8K1�/P�e3u�ʻ��`�J�/:����JO��� g�>V�D��ޫ��qI`���!+�L�V�G�=�w�W���j��o���9B��ldy?/��ڰ�Ֆ��iH�7�zN�7,���:�-b����.����s_�U����/5`�7S0�`꧳U�Cϐ�x�sҝ���ए�p�X���Z�Ar��1�7MF��j-�Ɇ2�1�����m:{�ȸ�(�5�=fIz)$<5����B,��Ѳ�%���}��d���#��e�m�uQ����H��ps�&"˽�2��S�]��,���N�(��v?�~���V�G�|[����#a���%d�)�"j`f�_=�צ!_�u�(E���*�-��*���@�IJsԗ����m�Z� �"p�����Q��iV:�?�`MH@���d��{t�M��q�6f;�K*��R� ��a�S[��ud	g��>�t��yE�Tʄ��/+夞�>vNoe�gz�e|W�r��{}��}��;��zTƗSZ�[��\0�_����e��ns�(N��K�t�-%�o������'���\���ajQ���b���D�2�޲C��˯j�A�c��
�ǭ�h�c��噴���Q���o�� '׼�����e4�X̗),��d�]>ߜ$�_FZlei�����Y��4��E?����h�*TK:�2�Cy�0���G�|Б�i<BKM�B��d ,���Wj%L�7,}Lλ�^T_����ư�ɯ�׋d��n�~mn��8���� ���ә��>�o�yN�fh9����I݄��#hM#NK��FZ�wv�LIIM!#;d������N���B�W��7=z����1Q��V{GRhva�=j��8�8��n�T�����@{���v8�3�,	���
���+�O��ѹضƺ�@���Ւ�-r���J�^��T�����0�GvnQYj癵%��2|�m�%�L]7:�_��&��(8���fn�ɪ1�
�eeE|#���D��a�O$�=��c�/�0.[�*��ef��䎯ً�Ą_kh9�B�b/c/0�r�T�@�ű����׹�`�J�0�3�1]��*{��Ϻ�@�Q��4Dr#2z��1;��>�"�@u(�w� �t�5��������2I���$Q�f��_���G�$Ѩ�ƛP�a��	�������rR>g��z�bS�	�z����	B��u��!�N�5N?%�$`)���7K�𣠦��Qޤ�S��V��F��!����&¶��m������C�udM327ZGE:�ܔ�Ӷ�l����e��U غj�f�Z�#�A��P9��������R��L�������J|V���Q`�:�g�m�Q���-���������mp��m88~�L��E3�1�Q�A=����4�X�Pj_a۬� ��?�N�r��k@'��W�7��g��.��'�Uhiv޻����\���#�9�}J|�$��u�v.��/�1�ͷ2"��V@gu��W@x9��E�./q{������_	n�p�{���u�heJf���ք�@�N�h�l���?Z
L:I�n�|���{Aé��͆YL\]/ꡒ�/�g�7�9�l����(�;`֧yr�[��v�����l�7pe8J�5��1#d�����	�ta�|�D�P8��t���'eb�l��*:���t<�I&M��nfx�H��^��������q�a-����(���b��`�uQ�P�2t%Ӆ \iOC�l̤l�����Cv���\ �k��%�Փ*�r<�-�&2꘻	��Y���Y�����K��a��h�/HtθH��Z�eu�6d�
F��|��}��b����ǚ.0��T���@E�}:6���<����rZ5���-X��)c��5��{%YA�/�֪���PK�`ǍLhJ��l7�} Y9�߂+A�������~�f�znlڍ�3|��py@����m�(i�*�T�-����I�&^R�!�5�AӹvA[�/o��ݫ�q9f�"�C=� �|vE���A����7�|\w�C�v������`s�Z,!�\�m���C�sߟH�_o��&c�������K\�~ 	��%���M��in?��~X5�1@)3�q��p���.T�l�\�����&����)��t����2�-�l�����q�$�&�;-��&��'���}=��M��ˉA�D�pҁ���Ȃ*�N��Z���T��M��`�������	B��Ң$�*��n�C��n� �i8.���e��s]���-���B��u��vw[�'قe}<�m(K�X/���
����ta;v�J����cƺ�����k}���i��].�m�P��]`���T���r�/�s�H������ �j�c����z�EJq�ob��#J�c/5G�F������Ȟ�N��B��.j�k��2��y�¼��@����D��㝑8
;��*�w	'�5Z���n�yI�z�O�����R�g�ٯ������9�r2�7v�*�,Q�*����BN"��3͟Af8C�|�"S-�IE>��⭪�}��'�{�ɷ	��;C��(;��%Jk�}��#��Lk�e�ux�u.�����bJs'���S��Դeײ�Z�I�
o.�Ruh\�(��#��m�c��U�f �L�fFE̀L�|NV�<��H���l$����,Y{���#��Zڪ��/Wc�zG�/.k�ހdz'�$��,M+��*e����V�l��t����v�����-=Z�@�v_T��9�0w�h�}E����d�!������!�n�D�3�~��R�	�b����S��r�U`�}鲺3>���k��g�ߡ%���n����I���/��r3�oe����s��S�W�Tq"�����*9=�*%���_f$�[:�âQ7� ���z.iwfT�* C��T�4�|�*��!���Ώ�;Z�z�\;`lo�ӷx�V�#�1�'�صL�%�\�]cG؈{�U�����6��f��(� ����5mX��>���By/�KdX|<���d�*1�M����0�:�U}��n_XCT�p�
{z��H�x1��Xf�ֿ�}�����|ܫ������ѹ2�3�gZ(�U�D6���0�����@�SW3��B���\�ǩw���g��S ԥ��~���(���R�e�n_�϶r��{�˲lL`�Q�$�N�щB>;��o��(
��I�FWI
�XӻD��Ȟ�a}���4M��]���Ǵ�ț%��-Ҕ����A�)�N��%�'�mUP �/r$�|��ա�~�G�)ld�-=u^\�Ij!�*�x��Ǣ�)��yW��O��:��1���d�!��x=�k�!��N���fp%U��~&�/�w�f�+z�ڞԆ�R�����oSa�eD� �D�L�[�ن�"h^��"��>bU7�q���y�����׌�׿�wu��E]""��l���#�D'�]��^�	���g����"*_:R�姛��ۊ��4�� =32ֆ���8�_����bǺŎ#d����k��U&���q����j2�?l�$�ڤG��?�?WM�[��6w�ܗw���oP�<'��8t�oZ0�Ǻ�%���n�xe��j�n��MR}ٮך����yp?jb5��OJ����	I�GM���*t+hM@Z�u��]�]��Sw�E�*-�ɦ����T�]TF��ծ�80�{kՇ�+�]�Z�7���Hç����,�y( 	�(IԸܻu�4I��
Y�y�F��1+����e�h4|y���U�P�������e��I#�Y�Ҝ:Z�Dk0�.ѱ;��s��9�/��b
٦,�T�������h�r����w�[8�'��lS��w�a��Z�ۀ�m��Gk��"�ET#�8:Wn��`M���C��X��-�SF�yM��A��]C��Μw�n��8S� ��~���@�-%�X�~>�|�Q�k��!�*Z�x�������a�/Zrw�b���p�8{+Hܔ����"�,�������`"�Z�����[[��A�8'�Z��%�4w�P���[x��?ZB������9NDR�w����P����OW�v��ϩ8�Wx$B�5(�C�E�#D�,���櫒=H�V�f�$���4�䬚-.�7��(�zA���N���5K|"�h�74���'ȏ�PE,�L(�ٝ��ޯO�+����<!8�H���R&���@$�[����C�P��/G��6���6`gp�R+���n�ak멊�s98�VI�&����4d���ٓQ�+ �q�}�z�-����zr��C��A�%�Az�d-b��E���y�"��+�����=��ZB�	>4h%p�!��$�IΌ��VdPa�/�	g�eO/B��'kZ�*�(�3��aL�����D�esG� �N���[�瞍����T���5��������D����2�]�.����x��������X&2�~Z�����d�'����M�QP���ڳsg���i�pM����ڰ�X/�5,��O��נ*����;��\�P�����:�A��zQBYl&1�p7�[�;q��md��2�{������d!��=�OGF�����٩�zk��y�v�M}�s5�4RnM��������T��=�?��;�߳���g�d1��ZR$)�])�2�B�#�h�_Q1�Z��e�9�O�2eU��'��M���bf�ʱ��}��]xK�F&u���s��B!9����JPA�Qc������>qpX�YHc�o�$�`���T٥�4�)4��{��5�O�b����Nn@���|����Q9��:��C�~X)[ܡv���1��v��c� *�Eô���_]ɳ������~��G���jtz+f�iĖ����lj���M-�3��?���w�p���g��tV�+ϧl��B���.�A�]i{���n���xq�Y�,e��1�j��*Za,����7׿������	q��w�����t�U'��qb
�$�o�c��A�[b�Զ������?w����z�JK��A���Xx�jo�D:в�
�� �ի:w��ju�;n��RU�<� �Xi ��6���
u��X�,�R������۩���nfy��-K�Ϻ���������:'L���<"�]���.�Ȫ[�oI=ʧ�3�9L�#���aw*?�X�YU2CF,pN��;�N=�������X_��8��즘y��,�@,.r�j���Kǖ���	��y��4���R4���a	T��� n�J�v%>�c�-�k��<���[�p9�jg�[))���<��SjD%�W�v�4�&s��B��8;3��qo� Y���F��B��%2q2j��!"f��`�鴕�95ȑ���x�ˎ^�&�˞t�j�]/��j)�Dg�fz'�`�s�if����F�7���ڤү,��q���Lp�yD!�;-���U�&m��I���M�`v�ˌ8��?�~
���pIC:5�պ��w���r���a�]�rcV���u/� �����)���>Z��Ğ(�x�|,˓H��°|��y�oR{�Wn�?ky�妾�I:�����i.�3x�b�̎�xp�d_,�U�l��Q��|K�Y�[y(�ܺA0��-Oym*.�t��0���Ǽ"5������Z��È԰��ɡ�6F�޸Ї!�f���n��\*I���!��7����~*�q��S�R��}����-�v�eY|�nb�Ny�d����G;����s�'5j$w��'���\�Nl��4~�1�5~=b5�W�Я�ju�Z���	�a�F�ʿ#��Y�֫[��l+HH�(Lƣ�b�%� �Ѫ�]�W �h3�@��0ɵX|۾���n3��L��3�#?q����@PG'���M��q1�q�Z�F��p��~��AE'�חzp�;�2��]�A,�ô�^�p��~^��)���5�]�$�j�N�����VA _6�hb��K�w��ɴ@K��T��W�_��0����z$�[Ήm�x���I涉�o��k"���K���@���N��km�G����e8��������w��U��.F�j �E�#+�^��.�
�\w Q��(@q�:��w�o���~��C���a����븡��s��İ5)⑂�Mn'dvN��u �ã��}䌬[zA��+����oL@3{�c|.�c����`���=�ʧ��*�|��"�(K��ܺ�x����I��r|��G��4�\�X"��g��b���:~���f`3�(������X���-v�a��Gb�ʙbá�l�g��h}�#f���w��<���չL����g�	V�+�	�����f^�p�V��T{����.Ζ����knēI�����gK�jG���6�����6�I�N@?Q��Q�Lwk�̥=wI�%��#ܹ�}��]c���Tb��(mV�8g
�k���kb�/���0z,-�{��pcR�$u�_�S��v��Z�-�<
�	yP��~���k<?�X�-;/W_��%�RǸy>K�s|���.֏%Q�W�࢞���h�X�YQ�cR�~L��U�%��8[���E�{�ſ�F<���8�T�99�**���$�5x���G&E���D\�g�r��֓S��k_�Mg�NKbE����. j�imA�FYA8���7=��;�OV%f�r�b�����B������� V�&����|\U��C4X9E�g��?���%�3�!I�]����8��{n���M�N����f�b���p_f�בTC?c���/���������)x!�!��73�m�ǔ ��(��˗Y(�!�7���i�|u&	�%'�:����e���c3���
W����-�	L~��~���/�{X�l=��qt�f�o���x4�p�n* RK��k(�I��3�\M�	��@�+��Z�����s�`W>�0m�$��
��O]D�se��L�}��a��-ܲ�o3ݬxs�C��݀.�ؓ�0G����QQP�fO���7|��U}I�w�;{���0�g�:�ϯ�l��P��9%t��+̢����ӲL;Iz�����|��.T��tcI�1IR�>1l������7������*b�s&$�I-��I���X�V���O>>>笠��W�ٞ�S*����|�?l�D��舷J��%X��e����[D���*��Mu��(�70�V ���*�n��2�B
Y����KT�禐JGбb3XwK��NdU�d�R. :k���$ld���ļU��8�4��[��.�	�&�0X5���d��ב��h� ��mH-�O�4��C=�oEF%9s\��w�W�Sv5{aCH�Ѽ������w��cfzG�Z�Q���O��x֦�b�4|[��x:�(jٍ������v�|�V%O��2�&�B ZHY]�F���%`��V�5�G�hwc����"רD���J��.� �7�+� �*:xhL�I
,��e7��1$�[8��l�k����q"��Eo1:o�&�:�ߎ�W�4* ��!���*k���Sȟ�KK�N��
�F��bH���:m�[øQ;6����xc*�R댵\��gY��t5W��� W��e5X�f��Ԇ�%����>%�z�'0@��c�!�~��`����~�l-���&��b�8ϛ�ǪuU@$�E�׌h��n��h`��iԝ�E�Y�lBe��ט'4�l�1��	���[�� ����͋W������_A��h9� ��;Ѿ���R'��	(6���� �[K��}�Ha�ugEa��1���:`�z5f�I{B�<P��N�jy�����t	m(Y�� n��n���D�_�OS�p˽~B��m�����_��xܨ�(��<��?9e��!�O��8���mU�-G2QzAH�O���#���b�Ѳg��>�=��A9R($�Xe�~]�sM�1���`����C���>{�5��a��?�����3}U& ��L��o�)jNr�`C���.D7k6���DŦ9n�bi���+vOgON"SyI��bt3����iZ��c=�-�_wy���u:1�M��_ë�O��*����{�X���v_
3,8�}�����B��ѹ�5��V6�ɽ�W2)5�Z5 �9�n�7��!�����0st��Ec��N�Ѯcc��p/���Wc��]�����9��i�7~�DBz�xU$6�ǝ���S��������F�n�}�qM$Mf�`�;;�D�h�������,��P�֘北G_�̥�h�R��A����K�T������#a��&t���X���'A�bކ�����y�Z���zW)��K�~��wS��K��,�_��q�遲{���ܜ�>��ea�4�A�����\ N�jT�!=�0�����j/A�B@q��E�Ӄ �����L�^�R�f�& ڴ���zX�Tݽ�au�l�9fJ�</v�8��4�����~�(�x��f?�'!�]�O���s��p3��u\��*8�O�Ư/<�h+���f&}�-�c�l��ߘ�6�;�v�+ʵX�9q��ZiG9&����.c^t�)���1�9��#
F���$�C%	�ך&4`E�$�_i��a?�;���|ۧ7�����b/k���� @/9�U�&�k��+��m���6K���>�J�GEy�7�����f���D�.JXE�t�@G�i��>�D����o|h����]=y���1��]��f�#R��b,=��T2��˅���,��枽��.1���m�`&�$J��M��@�7'eF�P�t&�$q��g^�ŊVy}0��W60{�&�i>ؖ���8?��[�6��4I"q"�1
�T?�u|���gѰ��sp}� &3:|�uY\�
�E���X��:f�Q��F����GR��1O?��A�7.l^=���,��K�"_��`�À 3Z6+�C�'[r�JH���I�nx���AC����w���OgNi �O���#��mq{/^=&�.��+���b��g��m`q=�W��]���đ����P�GnL�S��7�����j�YTc��e-]'˺��T$8!���[�- ����QY�a��y��C�����'y�"tl��0�A�P"�Ζ^��fһ��9rv(��q ��g���a��o��!^y��-"����A�:v��N���91;�b�?�l�Y�M�)���e�eR�6t5���e������g�D�q��=2ި���CwY��~�/K�A_�hH���"p�pj@��j/�%T>�U�ŏ�X�S��j�?�#߁^�a�D�_��Ǥh�^��g@�����y�g����BKh��m�tp��p���r���E��L��cO@�:%�^=�ʹ�`J�y�&pc&B�վeoBj�tHR�"��r'�IZ9�5A��G�̀�g���9㐃�Tlg�A=W�ZmD���� |��F��Lm�WN;�i�8�S'�����U˽�s��/w���+��	�|P�:�k��A����J�j�93�b�,���A|۞ )���C����l����XL���!�&>���e�t8kkz�j�  ;��r8�x�]���$��t$�1�w���x�dݵ,Ce�Uj��O����PC��	Dr$ɡVK��ñ�#v�@�o.*e%<[͵�cGYq����q��zyb�]^��n�	�~dX͗�����kګ��Nj���P�Ϋ}M����u�+&.��>wHKE�5�����-�z�MV�t}s1�wӨ:B�����3�&��}��ܬ�8�0
���`d��4�̯���x�\L�}<kчj5���?V�:^�������-����c�A��-��t�$}�yQٴ��M<}�����>Z�H�?���&�>���guRL��q'��}����7'�m�2�Nu��C6��JX<�Ҽ�-[�U��N'��o�p1�0�ZJ�}�i�+�ټ����<ԇ�+���J��n�\�M5{}���������qT�{�VG�K�~p�~���:D�l��Q^� ��D@�B���kۄ��O
�O��h��&V���0� WCN4�aYQL��Cd�,�	^k.e.q:!%���8X�7D�j$�c�&�P��4!s�����{p��"M�/���Cj7�|���xt�}��n����N*�߾y�~(�Cf�S�-O�@�����a֙�&3SW5\�O@Y��ɂo�;<ګ�Np0�G*��B����yW��S<w_M2�§�;�)��1C�d��s�qF�faa�V�h�n���BE c>����
��\�
92�M�Q}��R�(!&
t���C�k.Z�/�H�["XX�	�tc�R����)P����9O��E�D��nM^���0a�����B`J���֫-(�՞p6�?>«<�`z�xp���/u�7�A���2�������I��QP���1+(U�~c��E�>(��]���/&�2]�W$���s�B��@o���2�����D��e���+��:Jo��S43�=�ȓSZ���#����N��Tԏ1����X���D��b6�{��u���~��$BHt�.hhW�{׉3$$>'am�����
���n�r(
:V�!��A�ҟ�Y����|�v]�3���o�'(3G���^<vAB�����t�C��8
 WN�/�3�L٥��[��܀�曖�ďw̡@E=���i3�	E"�2�NFi��+�Zr����\ߌֵ+<-�N.y�ڱq4C�����x��(#ۖ�u�p
�'+(O!�{X�>
��I2c�|���ېON �fH�)[�WD����WPH���@�_Ʊ��e�U�&���)�%�]����J?�_J%0�D(��=		��wB9X��5aܴ��y-E1A|�X�q�y������ܲ.��lSh��� �aT��1`���C".����[V:x����KG��Q���é;�f��N�B8��x!��7�(m��/[0����!"���C�6}�Jucwa���h�΍�|Nf���]%��߬O3��L��{.��������ŕ����uz���R�����ƛ���A����E�Ӄ�W=s�T\?�D�C&$/ىN���Ơ�#�=fK`�!���ݳ�D���_�]lIu (đr�h`L,�8n��)��#G)�_��=�)�e�ٝ��� 垼�.<WS6��k����p*���3��+�P��̌��?!�����?������<G}0ҷU����%p/�5��W��q}��>h诠<�[����gP�Z��2xㄢ�F��"/tn&�}a�����Ā�KF�B�#m<�+_���0;��'��w���%z��nŤy�Gz��u�LgQ�(�%R0���t#��x��y���#�6�c�|+�ȿ^U��7��R���\2(���j'(վ�Ƨ�]�ū��UG6�E�K�	`�<�'G�t�UE�׸	�!���a"�R��Ȕ�Ŵ���*0ʶ��n�L�u)-ݾ��ѣ�)�嶤u�}��߭�n~;�*sXk0�F�ľ��5tSш~xA$����^�	Ň�Q3X�� ��i�繨i8�?U��ֻ�
���[B�b�,>�
�W�Y�f�9�QM��Ȱ+ы�x���6�'X��C4�&��j��3�+�9ж@q�dA�-�����D�ugki*� םG"xϓAqKȈ�Dv����>U�exg�@�S�eP����۱�i,��w��Q7D<�@U>�޽J�2���w�5��b,��x+ĺ����L�U�+�8��5;x�}���5j�a�n���}b��:o6���X��R,q���ّ������[;�>����+7�2�j. ����p�`{�^�W�ߊC.��n.�zQHd�F�18,���N���e]08�c� j�	1w�p�j>���ToUĔ�El�#�OٳK�߬�}]��Ц 	�ceR�W��w���5�C��@�'�?����a����T����{����[q�7γA�����A�G��v����.z9�3h�9�T9X{}��ƕ�iA�s8[�ܽ�*e<��q������ �+	d�Q/4��؇χ([R^W~�E��M�������D�A}�p������d�����=��]]�l�E��Z��sa	�����WI��ҟ����f�#?S7�b�7�X	6�l�'�t�%�}��=����q�P�����Tv+��^nl(�M�����0n��ˁ�s������K��pc����9j�u̡+ͫ�0+����F��r75��O�7t�;�8���l��F	>��:\�2����:������ T��<h%�������L�������A��^�Y�V�.3�N�>���ޟ&%�����6�ҳ�h��J[	�����z�h>�̅�J��kӸ�(�uY�4���<�/8mӿy����wc�M�A�-��g�&��;y]�b��e�ى�۪,�pN�B�~�xU7�&'8�ll�G0���*j�9BHKa6Rgf���W��}�e��T�#�<B=4�~�@���%��.D ��O�%��B�MYt.���Y!M�ʬ��"_<J�=���f����{��!<vgG��bw���-���S7|���ۋ��aN*���En���TLy��s�8A���;�?�^b�Zz�q��'��p��}�_���z$`Ј7���uU���1�6ATb�,� �X\g~
�EMŬw�킵�7Ԟ��W�~�B<i��Q�UPCX5� e���SK�O�I�]��#�؃4lI.b$�������-�`}�A!V@��#60q���}eG��	v�6�	�y��.��
g��Fg,pb�N�Y�J�������2畜z��D��DغF^�D���v7u��[�ضC����z���c�l]���i 欗W2�m�V��́y}}co�����23�A�*���t
3�&3�������E�2^dH+�O���]]/q!�i���6b��'G�K�Ms���iJ�@�-���ߕ��ˌn�k�كkU������rTl�w.�����_5i3:C47~�+�����
�R!�Sܞm-I������#v/��n��;�PX-g�}Ӽ����E��P��\ÇE��)����`i��DLcכy2#��h����:W,�%u��3anndЋI��r���3nٟ6��Y���S�[���e��,��*~p⨖�(�l�����o�� *�kN�J�"[F�����'xo������`��m��A�=@�א5�	%ͭP���Q���B=	�\����K�d�m��Y�)��?���3i���6�.�~sx3���@=��!S���2���i�K��q�2�5����V���o=kU��_?��8U\�qS~�%V�bP��Χ����E��H
�y�|�(�\F1��)֞�>�2���\g8�d_C���TZ�P�d��XJ-��������_ɵ~�,/O&I���o)�D2�aZY��9���1(�S�����]=Ll�"�?a�}�|�f�MÙ��hf���|Y�gv��X��(�������H-�"Ou���$���vu����42 H�t�fVVG4|���50z���mHR��+W����-X ·���1�p|ܕ�|ĤG�>Ѽ�EF4&c%��ǫ7/�+�#�+���j�㇂!��m�SԄ��]��1�ɻ���͋u+�T�r@}4+��9�UF-ɋ>9�\�� �vX�h��M\砯��rvR=Z`8�8�SW6uӂy����σ��Ԁ��"�.ĳ�Y%M>�ל����<؅�����JK�{��) �N���A0�ˮ�U����N\��Hd�ں֟���b��47D��c�z#��?���঎?3�Ҿ}!9�Ϗ�
�W�n�8QA���).@�5���a�W��{렂hO�ʳW�f≔V�)w��F�Y���"��q�����j��7��k$�s��<�0	|Q�y��[��`���9q��yX�Ez��mȂGy��a���"��d>��mkR����/�x��	c���ü�hˉ���Z���Җ�m�j�V��!(~�e'�����{��W�o�|aAɒ<8��Ed� �j�G��6�j�d����5d�tC� �]�9����'���L54a<���\�vba�5��랒��s'�:F�^sz'
��s�fM�|×���JAĔ�YbǑ�y�6�V����zB�
{ꙑc�tFIO@*���!�*-f-�=�	�}R<BžQ=HA1��<��)yT)��j�gR���4��r��Y��`7��T�x��:d��W�onh��ᨨ(��.!��Dć@J���OD[؆�a�TE��8��F�W�V�f�����r:���-��/��-�J�U���~���ī\�wr��:�r�~��T��!�Ѕt��HX������H�)�d�P?�B=J�݌u!;�H]��B�/�Y��C�}�.t7�혁���jg��>@�0bn���8겝<Jz��4����ӊ��T�Q�
4`^;/#�O7��?	��h*.���4�qm��g��*2:�|�,7j S�x���x w��N��Ě����x*�^��4�<|�����E(2&2Z��9�)B*|M�?u	2r�C5W��1�w�]���� gH���عiRdM�[@ϡ�8V���=ޟdW�ڐ�go{����r�^���jY�6��A��Kþ ������m�I���1�Xy����'ȥ���E�����H� �ȅւ�B�~Bnc�)��ʉ��Y���5U�
�������^昄���7�5��#�V*�l��Z�G-�J�бJ��:�ܙ�l����φLb{9qsD��-%�e��o�`UF"P5a���<{ʕ!��˸#4��~����<_�Q��(#	b�X&SMAx�q`��vC�C�lw�X�\h�6;�&�}e��+��'��>��ӗ�=44�ՉL ku`0��$%q�
�����r]��e�%��k��-�q�IMW3�����2q���I���xmC�B��0����e�P�7���n0v�~S2�	�k���\��'��ZȎ&�)������)��*��W�d�5�r�BN����(�Ũ�eÿ//�<�v^t	�z�67P��h3���!���).V�R��2]��e�� .�,Ӵ���ܗ�s��~C����ɭ���.�x��U.�I↷����~'�ҋ:�lC�'QT�7�^�<�rh�n/�Ӎ��@�m�*�?�W�I��*(�5�A�^Q�]��1Uu������w�U�DvI����.���@����!ǣ�{�U�q��OTL����w�QDrΕ��V�ߘ5^GőD�
�{�h�	I�Ѳ�lé���ڗ��4���}i>��Y�h��?�.z���cl�8E�C�a�d6+ {��@��C�A�N��B�X3#b��_(�Dd1�4��ָ�SY�C�e
	+{{G����ݧP�Ze��R�}P��Vi�}CRa��9@��ʜ��.Z����O�E�O�>���^�	��4_a"��CC�\�J��߲�߻�ka�b!̈́M�v ����v���Bp|������̇/e(�=ٹ/,d躍���6I��-]e�$��0�}������kڢS��R@Q����#�S�x���f1x}1��B���pH�r~�*�W�B_ZIK��`�ʝnHR� nr��ˠ�G�q�T;��.FD*��݋<В�cU�ӈ��p���s,p5v�ж��k����̾j�E��~�L��[H}[���M6����j����E��fi����4e���g��J�+JG�Ұ��{�f�VQ�Mƪ��7�=��[��kz 0�5������b<���w��^���:m�Ȍ�lI�;�J�مˣ.����"��L�VhJ�O~�-H���ˤ�	����k��vB:��v0��ͼq�>Y ���s)mte"��k��Pџ.(���ܧL`��H�u�bDn����z�'^Ԕ,���V���!���gG �-�����T��%��A����J�1*o�.禂����晻	�e�Zz%�x���Y���~�?�.�����a�/u�jyV�>^(�,ƻ]ġ]0*f�ɝΡ�>��|f�&����i���e,�5�'ť�|���=��wQ�G%9���^p9�B7$�GhÀ���V&Rc���X��P��ɾV��!55�4�h�UL�D��'�x훳�6Q�n��������=���"@"�A��%s+Y؅i}�j'���WiLÖ,݃S�6��u>�Bb�7=U��х!+�m�!˞@��k��!V�*c�	�+ķ!����k�q)&Q�����m�"�)��Qٱ`,(@�(����D�]��QI�|H@I|�~|���d��I9c,:��ƹ�৐%�R����p)_�����rЀ~8�S������s���H1����5R�6>29��W?0��,׮�J�

���r@q[6��L�F&P�ԡyӕ�V)K�V	8��<P��L�-V��|I!�O���������,e�Y43�Y�|��⫱ �n������8�s7=��?**šrp��32~V��Oh\�2z'�>hg�jl�J��Ke6G����6}�R�2�i~-V��y#�;� �'��p��)��*�$E��[�����C'��-�ؼ2y.l��
6M��છb��z'ib1
���g ������VRg��⾾��CB��s���U�&я�t������/��A�� MD����j�B˥!5p}���&`("Z�\4��"��Z�νK�('�֪�"�X,�j����`x���|Zڅt���=�T�lT	ߺ�g@�/��>��3�� ��]���3NfZf��������טO-g6�7~��V�Q����F�JH���?����t�E��#w�[�H�i!�^��`;�#С#nV��&�-�\Pr�0}��*�ƁE]���}���"���5_��� �M�$��/�(z	�O�i"C����|S���h�*P���]�7w�+fM�5���R����ttF�%�)�*�5��'C�M����>�8��laǑS�Ŭ�11Xwq��!�n�g�oס�|�|)�(�}j�뮿��g���N��U�%qSGo]!Vla�6�:p��Se��%4�R�J�EK}O��3�:ƽ����]~?A?�w�,bǺj'"%�3�V�wE�� ��On�8~S�B�����ߩ���D4J`<���	,�O�R�}EO8C_�T	U��^�{{7�Oi��u�@P9Q�T����Rhgc�%��#���	�)���e�ǊF+�{l�M����tV��b]�Y�k��3_�H��6|(ʒ�Z���>��S��c�e,$tD���HU�r얻@u�����\�DY�0
�5���j��{� @���n�OZ�8BeV���S�����a5?V��&w�ߒ7��ߴ��q�?p�����b��qG���욄`�U�7_���X��\o�ZJ:�]-��0�7�#��Ҏs�������[�BL�38���B4��	��I��%y�����da/�S
HMl��ӡ1�oX���ю�F!����E�Z�5|D������� �4Ub��9#@�+��}��e�HU3YXd>yeQ�)����2J�� r�t���df_�_�Tt܍��&�
7z��Cs	l�}e#1H�����dd��^��@�����m	��sIqn�WAa��G�4!
��:�`�ߣE������*ӳ	}ȁ	M����>�ϙS�
c�ēqɒ���ySQ?!z��l���!
�]����:�fCſ��C��{z�>g�YFe1����o\m��|��b�\�5�I�ߝ��2��ǚQ�*S'9��i���4sFK�Ԛ͟-�N�te�E":X���J"��[�-��b�
��$9@ ��d����/1��*�p�^N���(�'����&fJ�٪��"Uh��$�y��<�Ptp(���J�N�L��ʶrR��C�/���4���{��PQ�O��-j��`�gI�!jA� G۷Ή�W6�N���*�N����}����ee���2U�z�������Y�♲>�y�9I�\ܚ�g��^M��
�Hp)V�XP��`\���M��ø�[k��{2��Y#�	�ϡ`�4�I�0����;�t���KJ��	K�g&��s�w�=Z����_a�jFΤ]�gH����%8
?��o��?���	w6�8�:$p�sR=�����>zL	���5g���ս'|�O5�ll��]<�+b�D铀�i$qi�!r�;���ⷡbVm��@8��C�4����+��'t�Q���]y|����G�+�I`{}O�A�/�J��ٴ���ځ\��;_`�ޔ��K�ȃZ|J�*u0�$���׺��o.2��W`n�A�7��� |��Qp.�s�kj�4f��G�\nJļ$��I�q�k�8��T��HJL/y	:x`������#J���|I<��4%Rz�lX�d�s�]��yϬ���뱈ܛd�/Q���p���^̒�K�����U��o��ۄ*�����p�(���(��1<MϮ�'�P(��D�_���KH��I��,����E�LA�{�aO���2;Dr+���-��6Q͜:-�3Hy�r� y�Ɠn(��C(�nǉWALf�$^�:��{��w��No8��M�S�p\���[$+wl�9�}~���zU�;~(fE!R�rZ{F�\����C4�C̯X6��ͱ��x���G��8X͂K���u��sU՟�!CFo��é�E�67j������O��<�Rي��O�������L��>