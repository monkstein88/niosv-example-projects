��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a���?�;��ȎɌ�K�-B���b��Ƚ�/'��{��> ��	^FV�X�;^iQ;
x��}3�X�R��/�b#�x��*�"xH���M���'NX�䕇�,�{��m�D�\�%ߥ�$�Lo�:htuR��$E$�! ,��gm�:6F��1%JC�� ���uwJH�I�"w�e����o}H�Qʿ@'�1��k�l�ÊF
�G1����4�c̓�u�c�E	�Ԙp�r�|�a���w�7j�n
�n	�	������b�Q�����x����!09�\.K�ݩ��Ǳ�.U��9{��b@ʠ��A{Y�� *�usMZM��0q��:mޢAЯ�)�+��I���5�=6���Y�S�e|Zǧ/��:�!&W�wg�� Y�}�$�[�	�b�~��Q�zZ�pOJ�B��ݳ�(r��PHj��@�y����-X	�v70��Y&�8e���ݐ�`�'�[, �������,��K@D/��8!�����@j�6��+ţ��yp�����qh���+�J^�J*j�X���d+�j�'F��l�5[z�!����dnAe�����%QCS �L40k��據 ���$�9aȣ��nw���yY��oܬI6�*��a�����8-��mqo�x�)�5)��Z}C�h�D.]�Ptr+w7���ь�R�$����G�׷�Lpe:�kS�h¤)� VR�(�O��)l1�b���⍙#=)q��Wz��˿���)���d��
�h�S(T����;/?���G��/ɗ��+nW����3��	�g,2o��Q�}m<ڡ1��nz�ǻ1�ڴy��D���Ծ�"�(�f�VY�s ڍ�yY�pՇ��d4�r��\2P�b!hk��4�N� �ڏcQy�]�M����� ��Emy�lE��>,作a��b�Ch��Ō8uϹ�#������2�L_jU\	�/n!B◻Mt��%��K� �8兂++�d6��U��i�Q`",Y|r���U���V����l�_׭�3�f~�l�_U�x��0�F���%�����?��v�G�,	:��!ܧ�Y�a�}2�168�;05���΢��8�7y�e!����s����*���T�� y�\��<��.���4�1O��z�6�m��N�<�W�����зvx"�z�2GVTs0�T�6I��{�6c�lXN�A����w�a�\Gd+�)yH��R��ee?�tW����yAC�?6�ek�4��~��_oG�CG�Γ����6����m��m�&�rc�$KS��*@�>����\'���(h"�Ɩy�P!�B�qm��󏂠�cV��V�&�Ӎ�v!<рP��`,�f�G
?��:Al�AH��S�G|9;)��vo�c*ۮ�>^�#�b�q�p�ݔ-��b^[S*�3Y����%�?���+@��uBr���0�����Q*�iD�ȅ֗t�[�ܐ�&�)��:�.!���)hk���Ǫ lۀ{����v&|�.��� O]���4=�H\��YF�?8�&Z����3��~^��]St�W�y��tv�F�O��A���^��(U}��2�f�ى�=_���5���s��P�VDJS-y\����w����ݣ�/���s56�S��mjʙZ{��H�z�񙨓�[WZ��Z�s��� ����!v��H>�"n�}�$t���������۶�/�'��?�4J�.�'
��O��� {>����P ��&�5c��#՝1�e��26�/�mL�ze��Va�M��R�k2?E3��/|ykhOrƯ�_6�o1�g���L/�6I窕 ��8@�x�]�
2*Dd����S�f܀̛�g�u�1�����3m�l��E�K�,��,`�-�P�I[@������wUk�~z:��`'R���E�N\��8��SdCu��݋�Σ�7���&�R�;M2 ���H#?8[���]tw{.�(����jL�O�xB]=p��+W�V]/���s��(/�f�S���fޣ�`��lҪd��JW��_��X�+n�}��rVvE
#�@'�1,_+{����	�h�������X�uy< "W����m�	{^�]o뵤�v�8B�%k���̇LWF�W<:ZD')�Dl�o5�)��I��<�[��y�n*^���u�$_W[�O5DH�P��y(���n�3�=q��4�?u}P�#�����MR*���wj`J��n��E�����W���7$	�r̚����w?�H� �?k��<��+��^��=�����5�OK����!_����+��a�3�.���>��_J���Ceޛz��P���][��}J����x���(}�`	�Sɯ$F�"�H���nkͥ�?N{�cE���P�mN�Ot�粸�iГ���ZQ"����D��D�x�Q6N=?��=�"){���aIћ���{��"�~�����G�ql0T��>ӕ�X!_seCa|)I�J�\�c� l�����^������E�07��Z$@V�"P;���J`W�z�I��.d��pl+�z9ف������d�+�z��BƝ��X��W�Y;����	95lP��D�?��bTs��Ù��1��)��ֲ՛��#��=i���ڈ���f�}7h�-�2r@�Q��?T�'yR�L���z����_��lt.�jT�#k�;��%��V9�bׅo��mX[�ݝ�.�v���c"�ÒM���:��ek��^�Y��i�&���.���̽l�c�<�1T�����I+�'%�/�x��R���Έe	�?X=���xR���v�3�_�5.��	}cˤ��L�IP���q���n�����`۳{����g�2/�U�"bo���Q��O��1��]Fk$��,�ƐoZl�����:��t1/���3:� �w<��:y6\��{�L�V�hCڕ�O������S�n�is���av`�c��e�KN�#��u�4��a�5.�As�^�fz�������/�B�<���{�F�t'���)����òS�A|W�չ�Y,����/'�WurS��+���'���Jx���^������r�d)X�3OF�A0�1-w�?�)�ja�Oi�;�$��0z�	��o�^<n�F���n$�#��ᦥǃ�;�GL��3L9_g���lF�]�&]����qj��
l���&�	1�ɻ���_��5ߏ�9�=.jO�%ldov�Ojgd߭i=rM=���7��-�X�pMK#�����4#}��B�H��q���/�>>���%���M���ϛiҏs�3z9���`���>0��פ���>z�c7��O҅������Fj$�(�c,�aU�=#��ms���՞�ٿ��ސ���#IV1
U�%�F2�#(�g�h��K��Oz�`�/�?T�w?R�/{@�O�Z�όl?!˱�-���hJ�����d� ��<�~N0���ݨ�p�{��P�������q ��w8ۀd3@���PG
�"\5���ē��_~��!��)l���Q��WC�͕{�R|�&�4�Z�`D��W]GC�0���T2֗�O%���}�Y9��wӥ��AiOeW����/�| �1)�;4HC"�?����g�Z�v@A�!�o����>��x�L\�w�+Jjb�o٭���׋m�>~ ���dy�Cwk�?ۻ�

H��W�
���N�K�-�Lp�����)>��<̋L��׻7?S��z/N"�v����x`��3="r槁��.%����&���-S�g��z7�Xв�2a��s�Pz�Q����]ч��!�^=6�}�M�����q'4��5G�p\��AQj�vA?WrFQ܍��G��\A13mdԥ�����%��Z��Ԝ�]��.��D�Ny�7�my0R��*�t���q� ���9[U��B�Μ��>����G{M�to5�"�wl���Q�	V����%C8��HsfĢɧ�jr��d�r� g��~p��y�߻Cb��"��8�8vG,���
�sH�o��"Ea��O<��Ã�S���))�&KM�t�U��P��Np�?.�O).�y�yƁ�C��������MfP�Y��	j���rD�Gtt��Jk�}�C�/�H�?��#C�G���GO/
����pM�/5�А�jݟ섷�?/���{1�ܶ����L���,D{��^A��.C~�^��%qJ����Zj����^��B���;/3aI%�g/�J�� ���7j;�
V�3Z�_��>A��S٩K�!!L6z��u��i��}����G.P�Ȼ��L����	��%q��T�ٗ<�[n
���ȠQjw�o�C����x<ѱ��T=�(����h]t��Y���&�z,��_�Ty��|���������-ѣ�����G����>�)Ua���0|T�b�6PfW!6�rLv��4�Eg��Ɂ[�tD������>�Ǣ��hEtV��gE:dJ�Q�G�,R��%`��<��ҼxBX�2!�����i��0���f�*O�C^'�����ςM��O3���˦��u��`���i�"�tTfZ�%ZBkN��2��[U���%A"M6�
�)�֎L��zk@zj�5�*
jz�X�5M3�m?�I;��N��(l[�'9?���]v��!�˱�#Oے�I8.��54w��N����ٯ}��6$w�&_�C5�Mi�JЯ��9I��>;������6�c9��E8�d���fƳ-KN9@^h�zb6^��*��&i2��0���� �nR~&f�4ui귢c	k*$�Ka�;�3݋���	ø�i��^�:��W< �Y��i�9�*G�Z�l;�f6�ă���VӀ0d�:��w�t��Eı����%�|�-�7�&��mKz���A� �qm �Ϗ�=B�_���YU��aE��
4�������w臨��>�A�髪���hKL�Fڼ�Dp�K�힧\��g/M��+h�Y�LU�7�5x.'P������&��!٨ؠ�2��ʶ��n�Ղ��/ǝc�b�+�ROǭ���:��x���t���n��;�9����j�/�.���I����l?!�\o��4�t�Y@����p�Һ�zK��T����3��z����ü���Z-7�L�lg������5�M�����h\�	<�+�O(�����m05Q�(�w��9,��t��8��H��/�
ƭMn��w�v��&3�`��%9/8��ҥ$��g��B4W���0�@�h⏴K�`��E�v�l%�eNhlO��� ��qg"S-���y�,���Ԙ���'�t��{{6�KG�h>�6��Ǵk���"8&-�ff�+�[�TE���4���e_���.jv���!��M��Rpz�]�h	_C�`J὾����w<M_���3=�GQ���x���J��dzc��{��B}�ҳ��|}��a�,e��eA#��ҩT�F@>���3�O�o�(s�����m��+6��VD�ى�G�C�,���v�>���7p�:�ۜ����6*3���HR��T}�GQ�R����y� ݶ����2@��iګ��>CR�o��"�$�����޵�����򧼅j����'g��z�W$~�>I>�A�P��%g�rIDٶ7r_��0��&�H�ֲ����n���Zw���Y�]G��;�$�4��[���6滚%w��R�3���ӯ������h�wҤ���w3\X���+[�-�����έ��'��^^b�8����\
K�r��P�׎^�h��骵�w)
��Ň�}�ɮIGd��u��Rg=���U�������W~0�`���d�N{��5Ą( V`����9RP�/WG�AG�-�U�ꓰ%��h�����g�9/�2�����������&K`Α��2���Ӿ�o7�o��(|��"w����W�ڷ
�� #���S2�����b�t�3�82d�KI�$�;�]�nn[�^���w�S����HP:XV��rπ�c0Z!�vo����K�u�<��fg�@Aq;W�8G�L��]�N�V�<���1)N��*.R� �i0����!���G�`i��1��v'D΄�𕧣#��0�"��B�!)��/k�i2�\�؟n�A���y����)j~������m�W���Ć���6�'I�'Y���������-3��;]Rs�_�����]o�e�ր���;6��C���`����u�[m��J#�IA��
q�~;���<Q>'2��P~�7�U(�1��z�~��5n�����.�,�A�V�^<4�����g9.���f���B��+57��5m�}@�w����֞���J���[�=)1�x�+�B��AG�Rp��Q=b�7sF��[�����`�om�?���T���Hqt}��8��ǘh/}��߷$�ZƊf\��o!<Ie�|͆�i�u�A����/��؎!����i��:�^�𷁘�[�����QȎ��; �;���{!7�}e�j��xi��T�5��]O	 Eò�:��gɤ��CN��a��W��y�x��T�VU���J�B	TՆ�5���M�H���s���V)d��r�)X����?�Wq�+)ާ�$�.~�h�e6�8�f�踵C˘�̴���ٻ��n�|���hY^2�˰S��۱��� z&d�a��Ŕ}Æ�����U����G?��]��z��C\�5~�9֯������y0��י�7����(R< kU����CβQc�MZ�D��7��8�?�R��͉���4��6]%4�f��UM	o�+��������X@���L2�X�<�l?�8�!Qa�׺}p#�����:�(���x�T�F.�E���*^����Y�bӶ�Z�����zkM�~�6��~��%�B0�
��|�%ivvmDd��[�����0�>��x��=�pjC�)��l^l8=�n�K�O�a��-[����"��WSy�n�����~���OL���LK����m�H��^���F��O"���oQ�tj�M��.�qk4�Z���`��nX:�����{A�
/�h*����ǣ	y_��*j->Ѓ��6?�05AG|s���#�H$�1�2W�S���ı�=(V51:j~W8yN{��e�ʹ��p�:3�`�����uԫ}gf�m�����"��W�#��	
�v��7��y£�rh�+��X�{��n ��r���?�tc6ׄt�y;=��C���5��0;�D��4t�wO����g׈-��2��#��y��5���טh�/l�\dEq��������]s�h���/�W���VD�����s�K�S�b ��w�(~�/��r;Q4�G^9,��t۷�������/&#�P.��|��|�~���H��4O^7�vGR�W�yv��*�t�1�q�$�Kx��fgt���e.�Z6����C��'�a�R�eZP99���$~h��.��ʊK�v� '�&����,�^��o7�N��]	�����/1q�w%�_��e���y�I���Ƴ�<>�V5�ܥ\%�I���Xקź�����}%qڇ��9^��L}=
�ڣ
g23
B���B�����,�hnC
W�m����������'+S��&�a@i��$�3v��n��Kබq���� ^#�\�����m�Bɑ]�n
7�#I{S��d��=����\:*���i�87�!0t�UDpc�9��7y�`�-t��J�kGV|?/{��?�_Pt9����K318��,��l�`[Y(�ذ�X{���Z	�Į����������NM!fP����~�Φ���YĪ�V'�󛄜��c�)l�E����������nT�`��� Z�Eq1���6}+t�ᙁ@Q�\�}d_r�%�c�����hf�M��	>ɾ��z�TIX�p�$��P@�����LW�к���:���	L��/�pC�]���粫]�#�y	ԕ�7��a��J��'ؘ4�9��!��_A@� =\�VƎS9�G�¿hC����T��C�u�3�]��s�Ik�~`����?a��a��L~J%�R�f���#�n6��`ab&)�hgx?�������V�)���n�`���7p@(02�.{x/�:����ᥫdt��a0��_�]�َ;���N~l�S�S��ʻ$l@Թ�n�(�"u�"����X�(��d�����u��P��4: �`s#�C�9�X�}�Jx��T8��tU�y=�b�ON �%w[�Up_�eH
Jxz݋Cɠ݆��џlȱ}��!Wx�K��ZS�#|%�6^g��C�(s�Nxc�S�6��;�z�<�v��'N�A�S�>����o7�ĎE�fvŶD*n�qy8�kY�͙�W����Pr�V�|E�c2r$C���D +�ŝ-O{��.{Rw�`�a�ƯCU�J��JL��m]������I4����
�eg��;0���\�?9��w��
�ԅ�)��m����F=$�L�8+M^��� �|��WsH��o^%I;��/���(���7���ڦ��WÌ��vOxg�<����:̶3��G vI�~���a���~����qȀ�fҋ�"]K�Wha�Uv��j���پd;����zP�؋�C!���r� �d���{�c��(]1���Z6R{@z�zG�*�n���w�9_�c,D�{~���u[S*?1c��G���0h:���~F�+aϽ���S!�ߜX-�gH׉�/��>7��Fx?��z���k��9�:�M��Rt��7�Q`Y{}���l�(^���\�\؜E��M�.�άU��xy�U�gwU��mM�V,]�Q�m�>�+�JRr� Z#�
ސ��xH9�*J-��(o=y>#f_�i��!}���	�A9e��!�S�P�~��[��	�+����/��P����2\
�z=R�X#/����