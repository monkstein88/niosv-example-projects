// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
olfbsX6sNfi/habU+j4BJgR9t6ktjlgAJ3tvXZftWy+DZB+wHxEblQU99mwa6CMRfOTcMYmgn1Xs
qXI/QXqmDbaJVtyDB4j13Iqy04ZBP2rW9i2qWQA8XjM39hQ3UngHB+NqFS1r7L3yqcIAsS8+ed/E
tuF5MemJib+yd50Kj5V6RCboEDsfNhi1ij1s8zV1lKTs8hr4S177EQqY3bKst54wbfh3dLlD3IrR
EyS/1qzsX3ks/aDrjH0Nd1sTU4ULNqP4iDqA5Rv1P2+KqjT94JniJIHFkwAaGh5OBbXyltXqDX8u
C/KtDD4uNmlbZSjmGv/rqhrcC3Qa7k4MeL7Qog==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7728)
5Hie9q0R0ISiA6OvQu/bP+nJtmiLe2axQF7xRGwtZR6x3FMI+3AUhWNnN8Ggz/J3ONrq0X/1XUf9
6ZzEoDFi3DkJPGo+KnEMITiIbU/WCG5cV1XDSRX0EM3+Yv5F9KxNtxgBpLGM/RZWP2z9RplPtMlf
7Wttc0e6tDQQm+oqBNZ8Uqu/LO3+lbv5H0bOXmMZXCnV4EF4TYy7P2fzVWtF/XaGutTE2Z10COrJ
+IEXvzQKodTWKMmLtnzqqKD7oGh/ZDdMqDipQV8/wf/AgC0mbxqWwUUVTonzxe2SiocZIqcVZxN6
h5GzwTlfIdB2JEfkeBIK7xh+HfL0UXWHFi9nrOZ8iO55Eu9B9Ey0JDp2Y6SRqShm3l1vgsJEm9Qm
OtlH5wQ4KtjHdprxPtmKfbMe5+QOfrpL670fJrDPMarRgdZ53Y/yEy9rIrzD6gtk64rquCZcm2x+
JV1gJAZD11XTcEEvmNTjw8dhBsv8YoQl/wRDiDg7EhTEmNbdsH9rktG8B4zBcohiiRJgSze2ySQH
5IEyyKotafdmwA/PlwQDRHfoEwL81eRXYN1Jvj5fKKXYVXjs/3pybUBsLgfIL3ZJXUbzERydkycm
pu4m59VlUlwZqiVDakgvYqGXeqPnygimcHub/4jDwlz3a/IzPxD9oVoWoUTQwZ3WrK1iRe28VP7Y
mTwbQOUR9rp5VdnHCarFYPlO5YjSWY7nCaCKmBYWM21nUyd4jfgyxAjITg0YFOU9EQM1ZZi4xex+
w0e9gYrGoxwVpW5jZuHm48nR0xGVwPvdd2L7cSL8OGw5FJpHVvbp9kVWOXyMHW8saxyZ2H3g7PeH
q5n5oGXvwVMaoHwiYTlMi3oYgI9jpAuXuD2kTIGQYpp0xL6hFhp0shNu6mq6P2iIfybeJLvQAQcK
yr4Iburzdxfknk8UO2oEAG/GT+b6m0daKI2m1w1Qe9p4M/8zyE1nw2h2YjhND02meMSPG5s42QBK
RZW1ZMDWSVGQsk6CLH0oGsx2Wi0WRA/gjvyiI2icXRfV0B5/3r2tH4Yx9HQY8wJSlgZ9W7siASE7
VxlHQc7kpQw1Jb46Lq/mPvq9anvqB2JSnmxvUitp31PYjjvXxTcBcVtHwP+ZBl9wGRWYwBp9JZuA
d53byQHOP8ELa/d6hRpI1kL41goO4xtsnfVHJ1aAsV8I5/4KcgEhvcgKDMiprXH0AJzvOvXY0twq
vpv6xMopqoWN7qcO0hoTKQRAE4aVqYe9lUD/OizhWmEZcqjoQwboZo1A0ijH78xrHyks7EQarIfi
2A/Npenc6eiqorUFxqUbhBwk+42Mf+Vrp7IBFyHyoK+Q/G8yHiWCIEF88PfCHqVhX8vD0YGOq/Zu
L63UNof4RX2BUEJ8HpIi+rWqHq3NZqlv7rCErg84R+8alGhIVhczqitRrcyHsmFlEk340yVF/zZi
Pogc+8zfo9Trxe48I5nuF+HrGEX8XVunMAHKpPHhVyzeqcpojPNkh5PubcuLn0rcMJ4+zUIuome4
xhFtpKLJC0cyzcpGN2zjGwHHUzu0HHC3kejuw3Yd4NPjh8CGbSZGKxNNRynAmg1k0qQqgDHjRw4M
GzShFGtcgF2ZEXFnX9NBdpF1dopXNJs75M/eQEvP2sR94g5mlDX+UBKT5z6g0N96hJfkqpQoedkL
Sw4Hz84XLeOwNpInGFAgG2+op1Nh2jF9lDgVO6PTztBHFrEMsFlerLutBiUM8lcaXxvPjSGaYfoF
0Px8pKyC2/PzOKKVL2K+TAoaJB3vOKWG9ohqqFHa6kXNqCzksBTacecrLLht9NXbS6pdVB/S+hmt
WH8QJH+tYz73JtSvefXf1REAQHALD+GWSNNg9zihpldr4Ntfc5/pAqS6pVMJwTFc+VKBJSW/jeo8
wL43aCdJwYo/VZzDfKhr7K6rkmO66xOsJ0rhhj4MbYbjT61aFnL4G+9il3S3fTplSDV7HxAPrQBB
s45qoxsMHq1szgr2uO9XqmbCsoACz7U3if72z4xyzHIODU3dbQRweUNaM6nBxeC3XrEhfjn3kezr
2E/l8tdz0fDYOBHiTzUtM4Wx2HB8MFhH4UZlx8+oGj89I78pwenX+tNVWO1tYFb4kKEQsThfNCk/
7Yyx8/1ihL9CbqNFABsXt63QJoVyYLh3FFTXiN0veuVqbjcGK/R2RmMPi2sgU8L8vBgKcVdGpLwu
CjAc58N7YieN4/hTU93UX5rdtVKJ2gzppvNG9hF5jgx6X1EGmBqHyN4SPzFECagwucNyjX4HdLzu
kbdqUFKs07UEFm4mr8A2M63435gxShWT7DjXrGg6VsgihT7XNTuiuCldHXOYoOfpie4W2EMGj/ry
Jz7Yb9t7cFt+6tz+2QbLnyEWV0O7rEZMxBUiK0y9sNTeCQo5xFFYe714xiHOanQi+WRWM4wi7aVF
F5r872OKAaMVxYkHRz2GGPFU1L3iSsUBSGEDNCtV5WAdJufPvKz1L8o/srUkSSlvVVmqpXXjUwkz
owyGY4UlnaHI4DwaiBgE0d4MscHcEhMaNsM1BHyayCL7FtbnMLhz2jMXAaiKj3K+FNpfQwVkP0u6
XqJNVtasPeHIR9F9alFxdt62SFoRId4r13uiUzBDKuuAFQtAbFJg3t1CoO9kGOeOQWM0wEfdBnPL
6e//+C1ppfvAEDC5mteP6E1f/K578TtmAJ6cQpP2O+AhzurPUrgW0zP7RfUsyHNX//jXvZb7KJXL
LIlK3TcEPIDQUIF9dSj9wYkXEqO1epTmGOXxZxMXZDWzjK0+AcObHaGj4brVYqGTQGljcdYyTWwd
q7uhCFlRm4Th30ijJ5KmfW6kWoSNx9jzVHKrJLkyd+a1r++0nueLK/43CMJaTrsYkZJAKXSwRHUw
lLmhpoZkjY1HxWdeHTh1mqT8JnzAmCVJT9U44XbatiNcsDH2/NaFPaqjgXAl5qED3CbzDrmwUt72
lLosdKzpifIXbpvWZkHa7Pn0CDiSVqgSJ3yIg8smW4scD2nLwnKbzhSY0H3sukAU3niU+6iHpvnI
pbPctFbjd/rjOg6ZU5cjV8V9HKumjOne4pfKk4q4L99EmDmdCjDpIZnpP3F3up6TN7y57c16EI5t
1BAahOCtau1mDGUj4YoEJnc24Lkzo+POLSSXilcW8DwyNckDoz5yOcpFygwKCO3MlSdRgq1kNyhS
80nPDaVvEwU5RW8nOp3ou29fOEmKHxZyyu6V5l638aDGqZaiTbbn4nASK4/twm/5mOodxiuhLx9P
LRMNxS2ZXMmO6I85j5CyQr2nFpW+b8+GGlLv8ShJb2yC/48uWXiErxhv87wthlBCiVOsaI7tCJ5I
sPbiIqom0OwyOcejQmnct/Iie+iIRi8/SrPGcBkNl2BnA6an2K4Cmn3ifKZpsybIEsSLFccd4atW
lYK1krlZ07n+RRtd7aRPpJ09W6I4k7AzsaXmBmi9SZTVf2w24n6NlAInFSoX6ib4SUK8Zkr9IqPY
L017dy7P0bwnCQb8MFCBszDPOFi+mpZk75rQoyZIwdxlJNSUi0/klIHcSSEFXC9xlC4QHskwYJSM
6D81ZHfQkL3gFm08NrJY7rbflhgJuebkLvbxh6VQm/VtVc8g8rB6LjZ0+yhBFFYYQ3D1sfm9Ohyo
q34HfjqnKJVolwh2BKblEr807R80Eeyy4GfJbGdPEO2VUOvtaOKr4t+DfFk8yBcRVsfiTrl0mhq2
+F7d0ILUCK6rRDfuX4ls7frA5R43UdUzxvP6lIweOX+YASDcr3xGIyU1zGiwflRapbTJEZrMVGX2
RZwFybXrluIDXqSHlFs4MF/XZWfggOwWU2sF8y1DBEeNqpPj0Bn5j5OGmC2sw1sVj+eDj5N97+kw
FADTsJgtH3O3msSLtZsbhAJh6dOy+E5bD4VUJF/nYVhcvKFq8myfpGTBMHt/ujAr3l7WyPptvrxe
NwffA9gCOh8mupalP9ZINkSzgABmJCWbRhiddDeeHAdu5aEEFRhfbUgyF4oEuGIW7gpk1UA3rtSJ
M3eFEDCmOysYC828MPNHm6gHTIjl7xP/rExDZoxklmdsXu6wUlWyQvBdKQumaqwZeNaSqsF2g/f9
TN1XVCBqY+/xnaLWsTPTK78vkjef8oPnvZubPm9ZXDEn5OLDsGoMi5x3ZC3Fscdh5zm23+RmM7Lo
MwfoKU9YAh0cUPdYM4FTGcc1V0uckkRxl+v2BdDXdYfPd8ICHSpVXLSiRAve5ZXTQulj7nLExidt
1Pu9polHE/5cpAXWnQ/Uz6MQCBukYI8DEEFi3AdtRs5Z6kJfu8IKlvvovJCNxllNlp88FHffgk0v
h802me6EGA3VwA9Nleuya8Fy1ZY9eKeUTykIree3Qz4mHHMCV90GBXtTDQulNWhRHpfNrv2dj6gy
f+ndDfgRfsRn239HXXNVMuOerUXkHzBitZ58RvfP9fyGAhsU9eTsHJVMHJbr876YXRmqo+MA+7cM
MOoSpFNkSA2HqH9eRnOHmzjielaAtjlBVqaxQszFffzieAIf88lYwCdm7K8apkyI4OuTvkqgtpyF
Wsy8IKY1yFdhmv0Gaq6wRoF7kJUEHqUGVWcT/8GPOo2eqRomAldpJs7jlSwRbadfQ/dq91FsvFhf
f3jg7aeICmy4mzBInH9vWpyYzXwbJe1FlgErmMO1IFrBqkBW+BD1jk0u5E4g4Zhqc+odZt3Xi24E
+RLhE/xx2tUvuDPtOZOaKjqGtlc2Uv9eNk2AR7ar8sMss909ps9mBz2kX0wBDWKIRpMbpl1DxcGl
/dPcPk36TQdCNm7eZ6UXq2WDRjtPqxdH8opFq0Y/GLActKzSua2ZebAgMhu4zW4f1QAUFrHfr1Z6
7cYTLMxbAidXLLGypXjKp9xlBvI1Ya76tV3tcBqVXiWSbjrVTQo8lo/03jOm0Y5jhzKY6nE3iyc7
XZBXJVJ81QzVHHU94PMLnxOPCIJnE5lAh75KiHBCn9JSyvNUKoCUfskXn9LrzTaV3AO3nXOt+//Z
Ixegi74PcFtEX014CVWsmmF7eRIGTD5FyqaLH+fdTZklgw3cFzzuzJFwwNrmo1NiCdESqw0M1rK2
safz7tSj2erOYiOG2jqA+1VG9hwaOWQ4MEAGsnvn7Ai15mO+tDE15UZvGmRNyj8j67Gkm8e+JleM
Jc77mz1Up6U9E4F1DAhC3iiIvfCanWT2K+DPdFCJVrshKezMsWYBCM+iFzawUm4LHh76VJD6DxLJ
YTEQbxstZGpUTg/U5lhT8gqyxgnQsQ7OKAcPYjImrssCCYbaFtRRPnAY8rxZNK0KtWDwKkdsajLM
b6+yG3hDvKFxyDQ9j7mxKA6bf04jaWxzcdfo+g5Vscp9hfw8+hKZ83AvWzx5lEki+QDvk6GNXEKS
juP0T9nVEeY7/OAtgDn7u2AbgWHTmT8SMOBu+be4ps9I7Wt0+xzOeA0/vMwkOU++0ehAAk6l/1+Y
djrBOfWXJJQ7TSdIYuual7copBh1twBh+pl6WyUVN+QhCwTUyOI2XgkwJVwIphirZR4rYCiXjJMr
1Y2vwZOpkgsMpjtqgZp0AkqWY3/ADAzCA9xo//0EW9nxT7oWguUKaxC0Lrb8+Az4aSDrGyfUR2Ce
/caAKMYs1HyBy4oi5b0Z1tU/ymUEE1YaSaekPIgzL+94s6FMVkv/Crs5Up71Zpc+3IRP/oecJrsY
60LaEVmD5RlWyrCIbTKBjKQophUy31JLrkLMG4t59jD09eP/Lbiy5Y2dBxCPfIrfkYs8/k75nq4C
XtV7kFn0kqhUTy9EpjPqgaEU0LjU2h7dp1HYTI8zar8iAGEq06/XmtEZTW1OiScMemiM0/jgRv0k
pljtY/x5auJuln+HvMdaFQANbHD9tM1lHbTzt8c3Ntp9gRME8Y9cqHYfWjqWB313u2az26E7bjEA
Z04EGSKX5EeUsbkCIyWmgnFmNHGwruUKJg77z4vnhREzIbmWM6v5o2HiDXenbUCM2LMLdIvVX4NT
EodL7L3wCjwLO7cd0FHBRDogzBGlvQikkOTU9ejDt7rPg1IUeTkcY/ztz6ekiU0HaI3hFxnVwhPS
LgUwI1PkTPINLC0w5bQ3Z0k7xGlvP51aAykUahO4ne4ngwDGVLs2/uNI5MXjyCI40SYc2K3NRLVE
Bwsmqywh0I4obhZ/Ss4B15hddjHeGM3lJJa8Z+aE8IAY3pHAnwziLP3n7LnDbWMLm2waygLm1mkH
Dn+2cCPal+AbX0JOudB6t4vy6JgwI29DExe9kzn23n7e7v5yoWUYZGU2YJ935MJ0+l7fpo6JSWeq
anZorsVqfIZ+CwnCGQiEZg2TrSIgsucEY6W19LeZpu6DDhnmAZIxIcVljH98bXodZ+NL+pXNTwHM
Q+XRw8e+8F/jvRn3q6KtstwamMrGptfvsI6PTyNQU8aFiu4OfFhug3yEMWo3rS1xHE87KeZjfZOC
RqyEgtD7mS0u5CA48Ms39mBLz7EWbq2b7QbjrxNCFu57m9Xpw0PvanvfjXUnW3TT1JqXnkZlJG97
CYU+LKdNrdQu5Gi9puka5FE1PUngSk8kPV00jJxDB4426FJT+/GWPsOUUFiyJs2U0pNHzQyRF6RT
HPT2gMUZmBbNCUoc9446NTZSXs0m8tN51cFeyNDgzXvuMAm5VQG9zqJ6YpfCg+lqL9giHgT5QXvH
gTAUl/VkCcIIxeXYEs9c0J/FjHM1ZXUe9A5x43R0tt3R8vLE5v8Sir+EqXWxF1YOMOXEWKZRFMXo
1EtJgkeSMUm6T+5h1GB9UDFBMEDI6SjAKwousVlzTZH5JDinlZ07yGtOesSDBHDDQwJJvH3rB+gz
U1UA2tZnkKq6RSiLu+eGA7HtM5Bs89nemGPqztRAcEwN7ZGT3XYd4k6Sv763mIlpwucQ99j6hfyB
5P+KPZRlpKREWl7RQUxTDKSrRnyCgnpzozIVXArkr9/EIqQZz0OsUIkH5m94cC8kN/07gH+AFyPP
pnc51klUxU2u7wjF0BrdVEJ5KAtR7LoSNGvTuJOsFqrDtJKmAYyrKtd6kqnnw7HUFylm3/oaHJUo
lcXBp+GkR5eIUdotjI63lP2S16FlC8m2EnHeBGqO7EJ0qnrLGNcoCOLZaBjQjRofB37QYBkOJLAC
y7NHTpRlTjTAY+5dNH9NPLlBCHHVT8VfrDMqC9irsO7F9i9W0FtlA3ALUoJ9AgTtBLeYp+guNHwO
6E3m8SIvWUCPwxCQcEWv1VHI/BKNFWF7QVM4/v/jujS7b47MVchv2K8ZXbYDnQcSOdHTijgrsCKe
ZJ12DDrj9DXiLiq/nQX5AJzm4yiuXbj8taKESmGFERH0/ntYbdLYGJVmhAQ9Rfrp+iBTaw66aW8v
mAX7gTLPDGCjLmyDcE9ixcpgP55VxuQn1s/KxwYMzY4edO+hi4lukovplsH7FzAQVlEtjmnMdUJE
q/LW7MhZcuK1qdnqw6H0IwdtoolJfSD/CR3khjcl+rDe0G/1U3uxONBbYk8H36k33RirilAvh0/1
/50yWL2IgKPi1WbrvSJZFHmyYz2xsXbIPwyU55YR0MLUDiTNK0lxYayQjr6iQn7CN3QkryTKEs5V
BE9COco+ouzIHadUH/Ta1eQU+69wGoMqS97EGV7jzQa4ECNJU8BHgz9vRsi2JEZvzb7D6hTF1NXU
SyTKyAlU/fwucy3GuawtltsTaCcndJaXkM/b8hFc0Au9dBXkWXlwUISzvyr8sIJ57zcJkPBDe/4M
VS0DFn+g6WU3g/ha2pzLl4b7TBhzPRcQtqqJHuwzMGqUdbLOcx6nd2Pud+ZO431gR6XSQ6wyobX0
2mkh67U5FzskvADuy0K33xYC5AFLgm7kH7MPK2KgT1l5JW1+LKHVJpEharN2EMZzbJUjBkVmB3HZ
MhnUR9iAssZcnZyG3SkpX3Y7Fk0e5eCXLt4MEN4XleBNgcfL2qx6I5P0aQWJZbyc0hWWfgKycOeA
iBVG0zeR+Su3jy/pn/MLm1XzeeFbZp/WDC/28Nx2U/T+5qNAj3O+VqaVte2mp0vuPCwEndb7z0nJ
6Ecgffl7rLWPKBN0N4XI4dS2R7IMkd61GubuLMbrTE3AiDpc2Ag6M3JhP5ECGcKzo2AGYNuUayVe
bJJUDD1GHroJODRjOwdTdfhCLFev0Q4djvDDhk3Jzbhisdiqz9zRskhw1eS8nkGlTuZilLDYg1m4
FPp9SwoH6p7rFwHDJyV60r4Z8sAmSBilmABEfMLTlhdRbX10rY2WP2oqAYO6t+UI8TYNkdEnAZ3/
Na3U5vtuWDfznSTszpkNsaSADMWgOTAdp/vnu1pdy+dYumw7lK8FRDrQw1Fv/CQ12YSvr6Y8y4YL
kosZYFpj3RJ6hC45X5kBotwgeW9GpmN6JFQ8aWrb3hqJz/gUUbrZ4kRIz8R78Q84L/r19E9hd3mx
XPANoDOADuF+QQGqgwuGgaEmO9j+bt2W6dLqNO9oxY19lX3mvxbFWuygcfJY5UqqFApoXkKoZ+7Y
DAfJ38posEJn6EC5ccRaTb8vDUrXY9pWcWQUpQtF4m+PgxcC5QNiTbfpopGA7uVtaINLzAoMzsIA
1R9uHxclPOONKsTd/GTz60iNyHeKTWCp3h9+47/Ev8SfxLh3e6h5MfNZM4NZuWe5PXMy/1Y9AbvY
aVhR27rsFDxLoZXcaqjd4Vjb/I+3C/2GgSKiXLtCO/Mj0eWcQ4VNMeCm9Ww9drP0p0fbe+/+0is2
FsU4Cmf4CTmFkrFq21TrOG7daH7D3NFU2o2jZqvh34QzAHwKedFH5qTFzqTcq4yEoqgjNdyraPJg
Jw2dklxqO5ASAW9ePB+b562iVk6XJaYoEV6QGYU2CcTQaS0vhTMwv06dOIfVYmU2IKXIHGd3gxt+
ZikyME/HfCdIV4RXG/szaV3pRi0LPMKM+Z35qeott9b8R6DTQQPPnTrSPYItem9H2+3Ejn0n5cLL
RkkNp/3eE6vtuhon2j2lTsw86yEAgaHLZ53XjMSPIeAarymXE7s/ppR0RuRvAjJ+vJse2kJFfeAJ
muVSs1ifmYRFVtnOhLs+R0ActM3D7GeQJQv5voEcbW7MR3GG7KUt1v5ONqvGnkSfGmu+AyEcwc5+
F3MnXtEX8uv1lkJIAESAdZgEFp9vpbsANiWyPHA//I3YVF1eOrajQ9OLpBniJekewfx9xYqj9wyP
Ng8RL7geeMAtAXBxXZijZHW3conr367I8nEAOPTPw2sywcKSqdNd3TPoQEDa0TWZPCDBannf0y9Q
bxmbw6JuKvleu3uQG8R9ZsGqrXCG/i/G8B3yiQVWnfenc0hJDXJC18xvGojAvlCPT0qv9WVnT4rG
Y9XebjA9ZPKqQRygLsoRldPv17gEisAD2X4lNehwhgbjjaiE064QYG0KQS/HQQWb7ZBtrpM3r4d9
Fsb/yGKYzlhZTsAb53VWQCOHkYL7c3A9H9KtSz8vLo70vVyzFmz0tbcP8cLRkX1I8okAGS6vW8Rv
Mc9ALKoJbY54apW7nkT9zbxC10DhLD4XYEO9LTp+CT4BRLS/5xHdQoA1Xcx90RjIpELr/co+1BNS
t6q0vi0ZG+a4GX7ZvfSUpG2KtXN8Z02XsnoPjTE+PTPk1Yu7SjtOY8GDPaUiaNFy4fptxKOMF1pt
Z0wB6ChA00UCAz/ULIdheDckTOZbYuJKWT8niGfQzIQmikmQks1V6skusrpt0lodFXC3RzsnsnFG
S1o08BPjMsXsXPzuHuv5Bi5OF66aFsxEAn7H8+z22Zm9k/yFi/T2ih2uHwxu5EtNEv3ZZR7Ody8a
LNaAlDVwDYxmfP0Gp7na/2z1/wHRJ/VQheNZsBl2pUvJHvQmzHJ/88beV0nqpZlaRv8BFVgqaVvH
Ow1bdoU5chWB46ZRYGRyAS1FnNGUFO0vATcX9Au/H+qkGM0Ye1MMNlJYSgfgPapjX/Fl4aacYQn2
cxa6USnix3Ub5Tm9VaE/fd5DVlDMBPc8kbFy1dloJGlmDrSZXElHLu71E+vhKMNxqc02tnECRy8o
9CBcmWGcqJAFODqc1A8NfxqtYvRlvvB4DBiteQg2k76p34/JtF/kT2t6ML9EB9ym5XhrNIsGdjJU
hpIOW6Fq4IkaBAKrvhC+IJntzCV5CPLU0Rw7e1am+WyhUcB/RMqrlOadujSeaUHeeavu0oNTRfv4
FCTW/6KDdu3071WSWOGwXpmciWnfAkg0lx6dJRFQN6hpBSRPKp4fYDX7WkuCgnQhFQr8wq7ASSN7
M9e0ua1kfzdeV1ccGsMSPxyEpud/cmXEwOzdLkouRiPA
`pragma protect end_protected
