// NIOSV_G_SOC.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module NIOSV_G_SOC (
		input  wire       altpll_clks_areset_conduit_export, // altpll_clks_areset_conduit.export
		output wire       altpll_clks_locked_conduit_export, // altpll_clks_locked_conduit.export
		input  wire       clock_bridge_in_clk_clk,           //        clock_bridge_in_clk.clk
		input  wire       gpi0_btn_externals_export,         //         gpi0_btn_externals.export
		input  wire [3:0] gpi1_dipsw_externals_export,       //       gpi1_dipsw_externals.export
		output wire [7:0] gpo2_ledg_externals_export,        //        gpo2_ledg_externals.export
		input  wire       reset_bridge_in_reset_n_reset_n,   //    reset_bridge_in_reset_n.reset_n
		input  wire       serial_uart_com_externals_rxd,     //  serial_uart_com_externals.rxd
		output wire       serial_uart_com_externals_txd      //                           .txd
	);

	wire         altpll_clks_c0_clk;                                                 // ALTPLL_CLKS:c0 -> [GPI0_BTN:clk, GPI1_DIPSW:clk, GPO2_LEDG:clk, JTAG_UART_COM:clk, NIOSV_G_CPU:clk, SERIAL_UART_COM:clk, SOC_SYS_ID:clock, irq_mapper:clk, irq_synchronizer:sender_clk, mm_interconnect_0:ALTPLL_CLKS_c0_clk, rst_controller_001:clk]
	wire         altpll_clks_c2_clk;                                                 // ALTPLL_CLKS:c2 -> [EPCS_FLASH_CONTROLLER_PROG:clk, irq_synchronizer:receiver_clk, mm_interconnect_0:ALTPLL_CLKS_c2_clk, rst_controller:clk]
	wire   [7:0] niosv_g_cpu_data_manager_arlen;                                     // NIOSV_G_CPU:data_manager_arlen -> mm_interconnect_0:NIOSV_G_CPU_data_manager_arlen
	wire   [3:0] niosv_g_cpu_data_manager_wstrb;                                     // NIOSV_G_CPU:data_manager_wstrb -> mm_interconnect_0:NIOSV_G_CPU_data_manager_wstrb
	wire         niosv_g_cpu_data_manager_wready;                                    // mm_interconnect_0:NIOSV_G_CPU_data_manager_wready -> NIOSV_G_CPU:data_manager_wready
	wire         niosv_g_cpu_data_manager_rready;                                    // NIOSV_G_CPU:data_manager_rready -> mm_interconnect_0:NIOSV_G_CPU_data_manager_rready
	wire   [7:0] niosv_g_cpu_data_manager_awlen;                                     // NIOSV_G_CPU:data_manager_awlen -> mm_interconnect_0:NIOSV_G_CPU_data_manager_awlen
	wire         niosv_g_cpu_data_manager_wvalid;                                    // NIOSV_G_CPU:data_manager_wvalid -> mm_interconnect_0:NIOSV_G_CPU_data_manager_wvalid
	wire  [31:0] niosv_g_cpu_data_manager_araddr;                                    // NIOSV_G_CPU:data_manager_araddr -> mm_interconnect_0:NIOSV_G_CPU_data_manager_araddr
	wire   [2:0] niosv_g_cpu_data_manager_arprot;                                    // NIOSV_G_CPU:data_manager_arprot -> mm_interconnect_0:NIOSV_G_CPU_data_manager_arprot
	wire   [2:0] niosv_g_cpu_data_manager_awprot;                                    // NIOSV_G_CPU:data_manager_awprot -> mm_interconnect_0:NIOSV_G_CPU_data_manager_awprot
	wire  [31:0] niosv_g_cpu_data_manager_wdata;                                     // NIOSV_G_CPU:data_manager_wdata -> mm_interconnect_0:NIOSV_G_CPU_data_manager_wdata
	wire         niosv_g_cpu_data_manager_arvalid;                                   // NIOSV_G_CPU:data_manager_arvalid -> mm_interconnect_0:NIOSV_G_CPU_data_manager_arvalid
	wire  [31:0] niosv_g_cpu_data_manager_awaddr;                                    // NIOSV_G_CPU:data_manager_awaddr -> mm_interconnect_0:NIOSV_G_CPU_data_manager_awaddr
	wire   [1:0] niosv_g_cpu_data_manager_bresp;                                     // mm_interconnect_0:NIOSV_G_CPU_data_manager_bresp -> NIOSV_G_CPU:data_manager_bresp
	wire         niosv_g_cpu_data_manager_arready;                                   // mm_interconnect_0:NIOSV_G_CPU_data_manager_arready -> NIOSV_G_CPU:data_manager_arready
	wire  [31:0] niosv_g_cpu_data_manager_rdata;                                     // mm_interconnect_0:NIOSV_G_CPU_data_manager_rdata -> NIOSV_G_CPU:data_manager_rdata
	wire         niosv_g_cpu_data_manager_awready;                                   // mm_interconnect_0:NIOSV_G_CPU_data_manager_awready -> NIOSV_G_CPU:data_manager_awready
	wire   [2:0] niosv_g_cpu_data_manager_arsize;                                    // NIOSV_G_CPU:data_manager_arsize -> mm_interconnect_0:NIOSV_G_CPU_data_manager_arsize
	wire         niosv_g_cpu_data_manager_bready;                                    // NIOSV_G_CPU:data_manager_bready -> mm_interconnect_0:NIOSV_G_CPU_data_manager_bready
	wire         niosv_g_cpu_data_manager_rlast;                                     // mm_interconnect_0:NIOSV_G_CPU_data_manager_rlast -> NIOSV_G_CPU:data_manager_rlast
	wire         niosv_g_cpu_data_manager_wlast;                                     // NIOSV_G_CPU:data_manager_wlast -> mm_interconnect_0:NIOSV_G_CPU_data_manager_wlast
	wire   [1:0] niosv_g_cpu_data_manager_rresp;                                     // mm_interconnect_0:NIOSV_G_CPU_data_manager_rresp -> NIOSV_G_CPU:data_manager_rresp
	wire         niosv_g_cpu_data_manager_bvalid;                                    // mm_interconnect_0:NIOSV_G_CPU_data_manager_bvalid -> NIOSV_G_CPU:data_manager_bvalid
	wire   [2:0] niosv_g_cpu_data_manager_awsize;                                    // NIOSV_G_CPU:data_manager_awsize -> mm_interconnect_0:NIOSV_G_CPU_data_manager_awsize
	wire         niosv_g_cpu_data_manager_awvalid;                                   // NIOSV_G_CPU:data_manager_awvalid -> mm_interconnect_0:NIOSV_G_CPU_data_manager_awvalid
	wire         niosv_g_cpu_data_manager_rvalid;                                    // mm_interconnect_0:NIOSV_G_CPU_data_manager_rvalid -> NIOSV_G_CPU:data_manager_rvalid
	wire   [1:0] niosv_g_cpu_instruction_manager_awburst;                            // NIOSV_G_CPU:instruction_manager_awburst -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_awburst
	wire   [7:0] niosv_g_cpu_instruction_manager_arlen;                              // NIOSV_G_CPU:instruction_manager_arlen -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_arlen
	wire   [3:0] niosv_g_cpu_instruction_manager_wstrb;                              // NIOSV_G_CPU:instruction_manager_wstrb -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_wstrb
	wire         niosv_g_cpu_instruction_manager_wready;                             // mm_interconnect_0:NIOSV_G_CPU_instruction_manager_wready -> NIOSV_G_CPU:instruction_manager_wready
	wire         niosv_g_cpu_instruction_manager_rready;                             // NIOSV_G_CPU:instruction_manager_rready -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_rready
	wire   [7:0] niosv_g_cpu_instruction_manager_awlen;                              // NIOSV_G_CPU:instruction_manager_awlen -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_awlen
	wire         niosv_g_cpu_instruction_manager_wvalid;                             // NIOSV_G_CPU:instruction_manager_wvalid -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_wvalid
	wire  [31:0] niosv_g_cpu_instruction_manager_araddr;                             // NIOSV_G_CPU:instruction_manager_araddr -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_araddr
	wire   [2:0] niosv_g_cpu_instruction_manager_arprot;                             // NIOSV_G_CPU:instruction_manager_arprot -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_arprot
	wire   [2:0] niosv_g_cpu_instruction_manager_awprot;                             // NIOSV_G_CPU:instruction_manager_awprot -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_awprot
	wire  [31:0] niosv_g_cpu_instruction_manager_wdata;                              // NIOSV_G_CPU:instruction_manager_wdata -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_wdata
	wire         niosv_g_cpu_instruction_manager_arvalid;                            // NIOSV_G_CPU:instruction_manager_arvalid -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_arvalid
	wire  [31:0] niosv_g_cpu_instruction_manager_awaddr;                             // NIOSV_G_CPU:instruction_manager_awaddr -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_awaddr
	wire   [1:0] niosv_g_cpu_instruction_manager_bresp;                              // mm_interconnect_0:NIOSV_G_CPU_instruction_manager_bresp -> NIOSV_G_CPU:instruction_manager_bresp
	wire         niosv_g_cpu_instruction_manager_arready;                            // mm_interconnect_0:NIOSV_G_CPU_instruction_manager_arready -> NIOSV_G_CPU:instruction_manager_arready
	wire  [31:0] niosv_g_cpu_instruction_manager_rdata;                              // mm_interconnect_0:NIOSV_G_CPU_instruction_manager_rdata -> NIOSV_G_CPU:instruction_manager_rdata
	wire         niosv_g_cpu_instruction_manager_awready;                            // mm_interconnect_0:NIOSV_G_CPU_instruction_manager_awready -> NIOSV_G_CPU:instruction_manager_awready
	wire   [1:0] niosv_g_cpu_instruction_manager_arburst;                            // NIOSV_G_CPU:instruction_manager_arburst -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_arburst
	wire   [2:0] niosv_g_cpu_instruction_manager_arsize;                             // NIOSV_G_CPU:instruction_manager_arsize -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_arsize
	wire         niosv_g_cpu_instruction_manager_bready;                             // NIOSV_G_CPU:instruction_manager_bready -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_bready
	wire         niosv_g_cpu_instruction_manager_rlast;                              // mm_interconnect_0:NIOSV_G_CPU_instruction_manager_rlast -> NIOSV_G_CPU:instruction_manager_rlast
	wire         niosv_g_cpu_instruction_manager_wlast;                              // NIOSV_G_CPU:instruction_manager_wlast -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_wlast
	wire   [1:0] niosv_g_cpu_instruction_manager_rresp;                              // mm_interconnect_0:NIOSV_G_CPU_instruction_manager_rresp -> NIOSV_G_CPU:instruction_manager_rresp
	wire         niosv_g_cpu_instruction_manager_bvalid;                             // mm_interconnect_0:NIOSV_G_CPU_instruction_manager_bvalid -> NIOSV_G_CPU:instruction_manager_bvalid
	wire   [2:0] niosv_g_cpu_instruction_manager_awsize;                             // NIOSV_G_CPU:instruction_manager_awsize -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_awsize
	wire         niosv_g_cpu_instruction_manager_awvalid;                            // NIOSV_G_CPU:instruction_manager_awvalid -> mm_interconnect_0:NIOSV_G_CPU_instruction_manager_awvalid
	wire         niosv_g_cpu_instruction_manager_rvalid;                             // mm_interconnect_0:NIOSV_G_CPU_instruction_manager_rvalid -> NIOSV_G_CPU:instruction_manager_rvalid
	wire         mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_chipselect;       // mm_interconnect_0:JTAG_UART_COM_avalon_jtag_slave_chipselect -> JTAG_UART_COM:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_readdata;         // JTAG_UART_COM:av_readdata -> mm_interconnect_0:JTAG_UART_COM_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_waitrequest;      // JTAG_UART_COM:av_waitrequest -> mm_interconnect_0:JTAG_UART_COM_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_address;          // mm_interconnect_0:JTAG_UART_COM_avalon_jtag_slave_address -> JTAG_UART_COM:av_address
	wire         mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_read;             // mm_interconnect_0:JTAG_UART_COM_avalon_jtag_slave_read -> JTAG_UART_COM:av_read_n
	wire         mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_write;            // mm_interconnect_0:JTAG_UART_COM_avalon_jtag_slave_write -> JTAG_UART_COM:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_writedata;        // mm_interconnect_0:JTAG_UART_COM_avalon_jtag_slave_writedata -> JTAG_UART_COM:av_writedata
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_prog_avl_csr_readdata;      // EPCS_FLASH_CONTROLLER_PROG:avl_csr_rddata -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_csr_readdata
	wire         mm_interconnect_0_epcs_flash_controller_prog_avl_csr_waitrequest;   // EPCS_FLASH_CONTROLLER_PROG:avl_csr_waitrequest -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_csr_waitrequest
	wire   [2:0] mm_interconnect_0_epcs_flash_controller_prog_avl_csr_address;       // mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_csr_address -> EPCS_FLASH_CONTROLLER_PROG:avl_csr_addr
	wire         mm_interconnect_0_epcs_flash_controller_prog_avl_csr_read;          // mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_csr_read -> EPCS_FLASH_CONTROLLER_PROG:avl_csr_read
	wire         mm_interconnect_0_epcs_flash_controller_prog_avl_csr_readdatavalid; // EPCS_FLASH_CONTROLLER_PROG:avl_csr_rddata_valid -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_csr_readdatavalid
	wire         mm_interconnect_0_epcs_flash_controller_prog_avl_csr_write;         // mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_csr_write -> EPCS_FLASH_CONTROLLER_PROG:avl_csr_write
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_prog_avl_csr_writedata;     // mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_csr_writedata -> EPCS_FLASH_CONTROLLER_PROG:avl_csr_wrdata
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_prog_avl_mem_readdata;      // EPCS_FLASH_CONTROLLER_PROG:avl_mem_rddata -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_mem_readdata
	wire         mm_interconnect_0_epcs_flash_controller_prog_avl_mem_waitrequest;   // EPCS_FLASH_CONTROLLER_PROG:avl_mem_waitrequest -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_mem_waitrequest
	wire  [20:0] mm_interconnect_0_epcs_flash_controller_prog_avl_mem_address;       // mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_mem_address -> EPCS_FLASH_CONTROLLER_PROG:avl_mem_addr
	wire         mm_interconnect_0_epcs_flash_controller_prog_avl_mem_read;          // mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_mem_read -> EPCS_FLASH_CONTROLLER_PROG:avl_mem_read
	wire   [3:0] mm_interconnect_0_epcs_flash_controller_prog_avl_mem_byteenable;    // mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_mem_byteenable -> EPCS_FLASH_CONTROLLER_PROG:avl_mem_byteenable
	wire         mm_interconnect_0_epcs_flash_controller_prog_avl_mem_readdatavalid; // EPCS_FLASH_CONTROLLER_PROG:avl_mem_rddata_valid -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_mem_readdatavalid
	wire         mm_interconnect_0_epcs_flash_controller_prog_avl_mem_write;         // mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_mem_write -> EPCS_FLASH_CONTROLLER_PROG:avl_mem_write
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_prog_avl_mem_writedata;     // mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_mem_writedata -> EPCS_FLASH_CONTROLLER_PROG:avl_mem_wrdata
	wire   [6:0] mm_interconnect_0_epcs_flash_controller_prog_avl_mem_burstcount;    // mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_avl_mem_burstcount -> EPCS_FLASH_CONTROLLER_PROG:avl_mem_burstcount
	wire  [31:0] mm_interconnect_0_soc_sys_id_control_slave_readdata;                // SOC_SYS_ID:readdata -> mm_interconnect_0:SOC_SYS_ID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_soc_sys_id_control_slave_address;                 // mm_interconnect_0:SOC_SYS_ID_control_slave_address -> SOC_SYS_ID:address
	wire  [12:0] mm_interconnect_0_niosv_g_cpu_data_tcs1_awaddr;                     // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_awaddr -> NIOSV_G_CPU:data_tcs1_awaddr
	wire   [1:0] mm_interconnect_0_niosv_g_cpu_data_tcs1_bresp;                      // NIOSV_G_CPU:data_tcs1_bresp -> mm_interconnect_0:NIOSV_G_CPU_data_tcs1_bresp
	wire         mm_interconnect_0_niosv_g_cpu_data_tcs1_arready;                    // NIOSV_G_CPU:data_tcs1_arready -> mm_interconnect_0:NIOSV_G_CPU_data_tcs1_arready
	wire  [31:0] mm_interconnect_0_niosv_g_cpu_data_tcs1_rdata;                      // NIOSV_G_CPU:data_tcs1_rdata -> mm_interconnect_0:NIOSV_G_CPU_data_tcs1_rdata
	wire   [3:0] mm_interconnect_0_niosv_g_cpu_data_tcs1_wstrb;                      // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_wstrb -> NIOSV_G_CPU:data_tcs1_wstrb
	wire         mm_interconnect_0_niosv_g_cpu_data_tcs1_wready;                     // NIOSV_G_CPU:data_tcs1_wready -> mm_interconnect_0:NIOSV_G_CPU_data_tcs1_wready
	wire         mm_interconnect_0_niosv_g_cpu_data_tcs1_awready;                    // NIOSV_G_CPU:data_tcs1_awready -> mm_interconnect_0:NIOSV_G_CPU_data_tcs1_awready
	wire         mm_interconnect_0_niosv_g_cpu_data_tcs1_rready;                     // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_rready -> NIOSV_G_CPU:data_tcs1_rready
	wire         mm_interconnect_0_niosv_g_cpu_data_tcs1_bready;                     // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_bready -> NIOSV_G_CPU:data_tcs1_bready
	wire         mm_interconnect_0_niosv_g_cpu_data_tcs1_wvalid;                     // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_wvalid -> NIOSV_G_CPU:data_tcs1_wvalid
	wire  [12:0] mm_interconnect_0_niosv_g_cpu_data_tcs1_araddr;                     // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_araddr -> NIOSV_G_CPU:data_tcs1_araddr
	wire   [2:0] mm_interconnect_0_niosv_g_cpu_data_tcs1_arprot;                     // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_arprot -> NIOSV_G_CPU:data_tcs1_arprot
	wire   [1:0] mm_interconnect_0_niosv_g_cpu_data_tcs1_rresp;                      // NIOSV_G_CPU:data_tcs1_rresp -> mm_interconnect_0:NIOSV_G_CPU_data_tcs1_rresp
	wire   [2:0] mm_interconnect_0_niosv_g_cpu_data_tcs1_awprot;                     // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_awprot -> NIOSV_G_CPU:data_tcs1_awprot
	wire  [31:0] mm_interconnect_0_niosv_g_cpu_data_tcs1_wdata;                      // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_wdata -> NIOSV_G_CPU:data_tcs1_wdata
	wire         mm_interconnect_0_niosv_g_cpu_data_tcs1_arvalid;                    // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_arvalid -> NIOSV_G_CPU:data_tcs1_arvalid
	wire         mm_interconnect_0_niosv_g_cpu_data_tcs1_bvalid;                     // NIOSV_G_CPU:data_tcs1_bvalid -> mm_interconnect_0:NIOSV_G_CPU_data_tcs1_bvalid
	wire         mm_interconnect_0_niosv_g_cpu_data_tcs1_awvalid;                    // mm_interconnect_0:NIOSV_G_CPU_data_tcs1_awvalid -> NIOSV_G_CPU:data_tcs1_awvalid
	wire         mm_interconnect_0_niosv_g_cpu_data_tcs1_rvalid;                     // NIOSV_G_CPU:data_tcs1_rvalid -> mm_interconnect_0:NIOSV_G_CPU_data_tcs1_rvalid
	wire  [31:0] mm_interconnect_0_niosv_g_cpu_dm_agent_readdata;                    // NIOSV_G_CPU:dm_agent_readdata -> mm_interconnect_0:NIOSV_G_CPU_dm_agent_readdata
	wire         mm_interconnect_0_niosv_g_cpu_dm_agent_waitrequest;                 // NIOSV_G_CPU:dm_agent_waitrequest -> mm_interconnect_0:NIOSV_G_CPU_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_niosv_g_cpu_dm_agent_address;                     // mm_interconnect_0:NIOSV_G_CPU_dm_agent_address -> NIOSV_G_CPU:dm_agent_address
	wire         mm_interconnect_0_niosv_g_cpu_dm_agent_read;                        // mm_interconnect_0:NIOSV_G_CPU_dm_agent_read -> NIOSV_G_CPU:dm_agent_read
	wire         mm_interconnect_0_niosv_g_cpu_dm_agent_readdatavalid;               // NIOSV_G_CPU:dm_agent_readdatavalid -> mm_interconnect_0:NIOSV_G_CPU_dm_agent_readdatavalid
	wire         mm_interconnect_0_niosv_g_cpu_dm_agent_write;                       // mm_interconnect_0:NIOSV_G_CPU_dm_agent_write -> NIOSV_G_CPU:dm_agent_write
	wire  [31:0] mm_interconnect_0_niosv_g_cpu_dm_agent_writedata;                   // mm_interconnect_0:NIOSV_G_CPU_dm_agent_writedata -> NIOSV_G_CPU:dm_agent_writedata
	wire  [14:0] mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awaddr;              // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_awaddr -> NIOSV_G_CPU:instruction_tcs1_awaddr
	wire   [1:0] mm_interconnect_0_niosv_g_cpu_instruction_tcs1_bresp;               // NIOSV_G_CPU:instruction_tcs1_bresp -> mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_bresp
	wire         mm_interconnect_0_niosv_g_cpu_instruction_tcs1_arready;             // NIOSV_G_CPU:instruction_tcs1_arready -> mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_arready
	wire  [31:0] mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rdata;               // NIOSV_G_CPU:instruction_tcs1_rdata -> mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_rdata
	wire   [3:0] mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wstrb;               // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_wstrb -> NIOSV_G_CPU:instruction_tcs1_wstrb
	wire         mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wready;              // NIOSV_G_CPU:instruction_tcs1_wready -> mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_wready
	wire         mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awready;             // NIOSV_G_CPU:instruction_tcs1_awready -> mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_awready
	wire         mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rready;              // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_rready -> NIOSV_G_CPU:instruction_tcs1_rready
	wire         mm_interconnect_0_niosv_g_cpu_instruction_tcs1_bready;              // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_bready -> NIOSV_G_CPU:instruction_tcs1_bready
	wire         mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wvalid;              // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_wvalid -> NIOSV_G_CPU:instruction_tcs1_wvalid
	wire  [14:0] mm_interconnect_0_niosv_g_cpu_instruction_tcs1_araddr;              // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_araddr -> NIOSV_G_CPU:instruction_tcs1_araddr
	wire   [2:0] mm_interconnect_0_niosv_g_cpu_instruction_tcs1_arprot;              // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_arprot -> NIOSV_G_CPU:instruction_tcs1_arprot
	wire   [1:0] mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rresp;               // NIOSV_G_CPU:instruction_tcs1_rresp -> mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_rresp
	wire   [2:0] mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awprot;              // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_awprot -> NIOSV_G_CPU:instruction_tcs1_awprot
	wire  [31:0] mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wdata;               // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_wdata -> NIOSV_G_CPU:instruction_tcs1_wdata
	wire         mm_interconnect_0_niosv_g_cpu_instruction_tcs1_arvalid;             // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_arvalid -> NIOSV_G_CPU:instruction_tcs1_arvalid
	wire         mm_interconnect_0_niosv_g_cpu_instruction_tcs1_bvalid;              // NIOSV_G_CPU:instruction_tcs1_bvalid -> mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_bvalid
	wire         mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awvalid;             // mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_awvalid -> NIOSV_G_CPU:instruction_tcs1_awvalid
	wire         mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rvalid;              // NIOSV_G_CPU:instruction_tcs1_rvalid -> mm_interconnect_0:NIOSV_G_CPU_instruction_tcs1_rvalid
	wire  [31:0] mm_interconnect_0_altpll_clks_pll_slave_readdata;                   // ALTPLL_CLKS:readdata -> mm_interconnect_0:ALTPLL_CLKS_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_clks_pll_slave_address;                    // mm_interconnect_0:ALTPLL_CLKS_pll_slave_address -> ALTPLL_CLKS:address
	wire         mm_interconnect_0_altpll_clks_pll_slave_read;                       // mm_interconnect_0:ALTPLL_CLKS_pll_slave_read -> ALTPLL_CLKS:read
	wire         mm_interconnect_0_altpll_clks_pll_slave_write;                      // mm_interconnect_0:ALTPLL_CLKS_pll_slave_write -> ALTPLL_CLKS:write
	wire  [31:0] mm_interconnect_0_altpll_clks_pll_slave_writedata;                  // mm_interconnect_0:ALTPLL_CLKS_pll_slave_writedata -> ALTPLL_CLKS:writedata
	wire         mm_interconnect_0_serial_uart_com_s1_chipselect;                    // mm_interconnect_0:SERIAL_UART_COM_s1_chipselect -> SERIAL_UART_COM:chipselect
	wire  [15:0] mm_interconnect_0_serial_uart_com_s1_readdata;                      // SERIAL_UART_COM:readdata -> mm_interconnect_0:SERIAL_UART_COM_s1_readdata
	wire   [2:0] mm_interconnect_0_serial_uart_com_s1_address;                       // mm_interconnect_0:SERIAL_UART_COM_s1_address -> SERIAL_UART_COM:address
	wire         mm_interconnect_0_serial_uart_com_s1_read;                          // mm_interconnect_0:SERIAL_UART_COM_s1_read -> SERIAL_UART_COM:read_n
	wire         mm_interconnect_0_serial_uart_com_s1_begintransfer;                 // mm_interconnect_0:SERIAL_UART_COM_s1_begintransfer -> SERIAL_UART_COM:begintransfer
	wire         mm_interconnect_0_serial_uart_com_s1_write;                         // mm_interconnect_0:SERIAL_UART_COM_s1_write -> SERIAL_UART_COM:write_n
	wire  [15:0] mm_interconnect_0_serial_uart_com_s1_writedata;                     // mm_interconnect_0:SERIAL_UART_COM_s1_writedata -> SERIAL_UART_COM:writedata
	wire         mm_interconnect_0_gpi0_btn_s1_chipselect;                           // mm_interconnect_0:GPI0_BTN_s1_chipselect -> GPI0_BTN:chipselect
	wire  [31:0] mm_interconnect_0_gpi0_btn_s1_readdata;                             // GPI0_BTN:readdata -> mm_interconnect_0:GPI0_BTN_s1_readdata
	wire   [1:0] mm_interconnect_0_gpi0_btn_s1_address;                              // mm_interconnect_0:GPI0_BTN_s1_address -> GPI0_BTN:address
	wire         mm_interconnect_0_gpi0_btn_s1_write;                                // mm_interconnect_0:GPI0_BTN_s1_write -> GPI0_BTN:write_n
	wire  [31:0] mm_interconnect_0_gpi0_btn_s1_writedata;                            // mm_interconnect_0:GPI0_BTN_s1_writedata -> GPI0_BTN:writedata
	wire         mm_interconnect_0_gpi1_dipsw_s1_chipselect;                         // mm_interconnect_0:GPI1_DIPSW_s1_chipselect -> GPI1_DIPSW:chipselect
	wire  [31:0] mm_interconnect_0_gpi1_dipsw_s1_readdata;                           // GPI1_DIPSW:readdata -> mm_interconnect_0:GPI1_DIPSW_s1_readdata
	wire   [1:0] mm_interconnect_0_gpi1_dipsw_s1_address;                            // mm_interconnect_0:GPI1_DIPSW_s1_address -> GPI1_DIPSW:address
	wire         mm_interconnect_0_gpi1_dipsw_s1_write;                              // mm_interconnect_0:GPI1_DIPSW_s1_write -> GPI1_DIPSW:write_n
	wire  [31:0] mm_interconnect_0_gpi1_dipsw_s1_writedata;                          // mm_interconnect_0:GPI1_DIPSW_s1_writedata -> GPI1_DIPSW:writedata
	wire         mm_interconnect_0_gpo2_ledg_s1_chipselect;                          // mm_interconnect_0:GPO2_LEDG_s1_chipselect -> GPO2_LEDG:chipselect
	wire  [31:0] mm_interconnect_0_gpo2_ledg_s1_readdata;                            // GPO2_LEDG:readdata -> mm_interconnect_0:GPO2_LEDG_s1_readdata
	wire   [2:0] mm_interconnect_0_gpo2_ledg_s1_address;                             // mm_interconnect_0:GPO2_LEDG_s1_address -> GPO2_LEDG:address
	wire         mm_interconnect_0_gpo2_ledg_s1_write;                               // mm_interconnect_0:GPO2_LEDG_s1_write -> GPO2_LEDG:write_n
	wire  [31:0] mm_interconnect_0_gpo2_ledg_s1_writedata;                           // mm_interconnect_0:GPO2_LEDG_s1_writedata -> GPO2_LEDG:writedata
	wire  [31:0] mm_interconnect_0_niosv_g_cpu_timer_sw_agent_readdata;              // NIOSV_G_CPU:timer_sw_agent_readdata -> mm_interconnect_0:NIOSV_G_CPU_timer_sw_agent_readdata
	wire         mm_interconnect_0_niosv_g_cpu_timer_sw_agent_waitrequest;           // NIOSV_G_CPU:timer_sw_agent_waitrequest -> mm_interconnect_0:NIOSV_G_CPU_timer_sw_agent_waitrequest
	wire   [5:0] mm_interconnect_0_niosv_g_cpu_timer_sw_agent_address;               // mm_interconnect_0:NIOSV_G_CPU_timer_sw_agent_address -> NIOSV_G_CPU:timer_sw_agent_address
	wire         mm_interconnect_0_niosv_g_cpu_timer_sw_agent_read;                  // mm_interconnect_0:NIOSV_G_CPU_timer_sw_agent_read -> NIOSV_G_CPU:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_niosv_g_cpu_timer_sw_agent_byteenable;            // mm_interconnect_0:NIOSV_G_CPU_timer_sw_agent_byteenable -> NIOSV_G_CPU:timer_sw_agent_byteenable
	wire         mm_interconnect_0_niosv_g_cpu_timer_sw_agent_readdatavalid;         // NIOSV_G_CPU:timer_sw_agent_readdatavalid -> mm_interconnect_0:NIOSV_G_CPU_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_niosv_g_cpu_timer_sw_agent_write;                 // mm_interconnect_0:NIOSV_G_CPU_timer_sw_agent_write -> NIOSV_G_CPU:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_niosv_g_cpu_timer_sw_agent_writedata;             // mm_interconnect_0:NIOSV_G_CPU_timer_sw_agent_writedata -> NIOSV_G_CPU:timer_sw_agent_writedata
	wire         irq_mapper_receiver1_irq;                                           // JTAG_UART_COM:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                           // SERIAL_UART_COM:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                           // GPI0_BTN:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                           // GPI1_DIPSW:irq -> irq_mapper:receiver4_irq
	wire  [15:0] niosv_g_cpu_platform_irq_rx_irq;                                    // irq_mapper:sender_irq -> NIOSV_G_CPU:platform_irq_rx_irq
	wire         irq_mapper_receiver0_irq;                                           // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                      // EPCS_FLASH_CONTROLLER_PROG:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [EPCS_FLASH_CONTROLLER_PROG:reset_n, irq_synchronizer:receiver_reset, mm_interconnect_0:EPCS_FLASH_CONTROLLER_PROG_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                 // rst_controller_001:reset_out -> [GPI0_BTN:reset_n, GPI1_DIPSW:reset_n, GPO2_LEDG:reset_n, JTAG_UART_COM:rst_n, NIOSV_G_CPU:reset_reset, SERIAL_UART_COM:reset_n, SOC_SYS_ID:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:NIOSV_G_CPU_reset_reset_bridge_in_reset_reset]

	NIOSV_G_SOC_ALTPLL_CLKS altpll_clks (
		.clk                (clock_bridge_in_clk_clk),                           //       inclk_interface.clk
		.reset              (~reset_bridge_in_reset_n_reset_n),                  // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_clks_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_clks_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_clks_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_clks_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_clks_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_clks_c0_clk),                                //                    c0.clk
		.c2                 (altpll_clks_c2_clk),                                //                    c2.clk
		.areset             (altpll_clks_areset_conduit_export),                 //        areset_conduit.export
		.locked             (altpll_clks_locked_conduit_export),                 //        locked_conduit.export
		.c1                 (),                                                  //            c1_conduit.export
		.scandone           (),                                                  //           (terminated)
		.scandataout        (),                                                  //           (terminated)
		.phasedone          (),                                                  //           (terminated)
		.phasecounterselect (4'b0000),                                           //           (terminated)
		.phaseupdown        (1'b0),                                              //           (terminated)
		.phasestep          (1'b0),                                              //           (terminated)
		.scanclk            (1'b0),                                              //           (terminated)
		.scanclkena         (1'b0),                                              //           (terminated)
		.scandata           (1'b0),                                              //           (terminated)
		.configupdate       (1'b0)                                               //           (terminated)
	);

	NIOSV_G_SOC_EPCS_FLASH_CONTROLLER_PROG #(
		.DEVICE_FAMILY     ("Cyclone IV E"),
		.ASI_WIDTH         (1),
		.CS_WIDTH          (1),
		.ADDR_WIDTH        (21),
		.ASMI_ADDR_WIDTH   (24),
		.ENABLE_4BYTE_ADDR (0),
		.CHIP_SELS         (1)
	) epcs_flash_controller_prog (
		.clk                  (altpll_clks_c2_clk),                                                 //       clock_sink.clk
		.reset_n              (~rst_controller_reset_out_reset),                                    //            reset.reset_n
		.avl_csr_read         (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_read),          //          avl_csr.read
		.avl_csr_waitrequest  (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_waitrequest),   //                 .waitrequest
		.avl_csr_write        (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_write),         //                 .write
		.avl_csr_addr         (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_address),       //                 .address
		.avl_csr_wrdata       (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_writedata),     //                 .writedata
		.avl_csr_rddata       (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_readdata),      //                 .readdata
		.avl_csr_rddata_valid (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_readdatavalid), //                 .readdatavalid
		.avl_mem_write        (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_write),         //          avl_mem.write
		.avl_mem_burstcount   (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_burstcount),    //                 .burstcount
		.avl_mem_waitrequest  (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_waitrequest),   //                 .waitrequest
		.avl_mem_read         (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_read),          //                 .read
		.avl_mem_addr         (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_address),       //                 .address
		.avl_mem_wrdata       (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_writedata),     //                 .writedata
		.avl_mem_rddata       (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_readdata),      //                 .readdata
		.avl_mem_rddata_valid (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_readdatavalid), //                 .readdatavalid
		.avl_mem_byteenable   (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_byteenable),    //                 .byteenable
		.irq                  (irq_synchronizer_receiver_irq)                                       // interrupt_sender.irq
	);

	NIOSV_G_SOC_GPI0_BTN gpi0_btn (
		.clk        (altpll_clks_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_gpi0_btn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpi0_btn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpi0_btn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpi0_btn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpi0_btn_s1_readdata),   //                    .readdata
		.in_port    (gpi0_btn_externals_export),                // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                  //                 irq.irq
	);

	NIOSV_G_SOC_GPI1_DIPSW gpi1_dipsw (
		.clk        (altpll_clks_c0_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_gpi1_dipsw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpi1_dipsw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpi1_dipsw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpi1_dipsw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpi1_dipsw_s1_readdata),   //                    .readdata
		.in_port    (gpi1_dipsw_externals_export),                // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                    //                 irq.irq
	);

	NIOSV_G_SOC_GPO2_LEDG gpo2_ledg (
		.clk        (altpll_clks_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_gpo2_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpo2_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpo2_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpo2_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpo2_ledg_s1_readdata),   //                    .readdata
		.out_port   (gpo2_ledg_externals_export)                 // external_connection.export
	);

	NIOSV_G_SOC_JTAG_UART_COM jtag_uart_com (
		.clk            (altpll_clks_c0_clk),                                            //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                       //               irq.irq
	);

	NIOSV_G_SOC_NIOSV_G_CPU niosv_g_cpu (
		.clk                          (altpll_clks_c0_clk),                                         //                 clk.clk
		.reset_reset                  (rst_controller_001_reset_out_reset),                         //               reset.reset
		.platform_irq_rx_irq          (niosv_g_cpu_platform_irq_rx_irq),                            //     platform_irq_rx.irq
		.instruction_manager_awaddr   (niosv_g_cpu_instruction_manager_awaddr),                     // instruction_manager.awaddr
		.instruction_manager_awsize   (niosv_g_cpu_instruction_manager_awsize),                     //                    .awsize
		.instruction_manager_awlen    (niosv_g_cpu_instruction_manager_awlen),                      //                    .awlen
		.instruction_manager_awprot   (niosv_g_cpu_instruction_manager_awprot),                     //                    .awprot
		.instruction_manager_awvalid  (niosv_g_cpu_instruction_manager_awvalid),                    //                    .awvalid
		.instruction_manager_awburst  (niosv_g_cpu_instruction_manager_awburst),                    //                    .awburst
		.instruction_manager_awready  (niosv_g_cpu_instruction_manager_awready),                    //                    .awready
		.instruction_manager_wdata    (niosv_g_cpu_instruction_manager_wdata),                      //                    .wdata
		.instruction_manager_wstrb    (niosv_g_cpu_instruction_manager_wstrb),                      //                    .wstrb
		.instruction_manager_wlast    (niosv_g_cpu_instruction_manager_wlast),                      //                    .wlast
		.instruction_manager_wvalid   (niosv_g_cpu_instruction_manager_wvalid),                     //                    .wvalid
		.instruction_manager_wready   (niosv_g_cpu_instruction_manager_wready),                     //                    .wready
		.instruction_manager_bresp    (niosv_g_cpu_instruction_manager_bresp),                      //                    .bresp
		.instruction_manager_bvalid   (niosv_g_cpu_instruction_manager_bvalid),                     //                    .bvalid
		.instruction_manager_bready   (niosv_g_cpu_instruction_manager_bready),                     //                    .bready
		.instruction_manager_araddr   (niosv_g_cpu_instruction_manager_araddr),                     //                    .araddr
		.instruction_manager_arsize   (niosv_g_cpu_instruction_manager_arsize),                     //                    .arsize
		.instruction_manager_arlen    (niosv_g_cpu_instruction_manager_arlen),                      //                    .arlen
		.instruction_manager_arprot   (niosv_g_cpu_instruction_manager_arprot),                     //                    .arprot
		.instruction_manager_arvalid  (niosv_g_cpu_instruction_manager_arvalid),                    //                    .arvalid
		.instruction_manager_arburst  (niosv_g_cpu_instruction_manager_arburst),                    //                    .arburst
		.instruction_manager_arready  (niosv_g_cpu_instruction_manager_arready),                    //                    .arready
		.instruction_manager_rdata    (niosv_g_cpu_instruction_manager_rdata),                      //                    .rdata
		.instruction_manager_rresp    (niosv_g_cpu_instruction_manager_rresp),                      //                    .rresp
		.instruction_manager_rvalid   (niosv_g_cpu_instruction_manager_rvalid),                     //                    .rvalid
		.instruction_manager_rready   (niosv_g_cpu_instruction_manager_rready),                     //                    .rready
		.instruction_manager_rlast    (niosv_g_cpu_instruction_manager_rlast),                      //                    .rlast
		.data_manager_awaddr          (niosv_g_cpu_data_manager_awaddr),                            //        data_manager.awaddr
		.data_manager_awsize          (niosv_g_cpu_data_manager_awsize),                            //                    .awsize
		.data_manager_awlen           (niosv_g_cpu_data_manager_awlen),                             //                    .awlen
		.data_manager_awprot          (niosv_g_cpu_data_manager_awprot),                            //                    .awprot
		.data_manager_awvalid         (niosv_g_cpu_data_manager_awvalid),                           //                    .awvalid
		.data_manager_awready         (niosv_g_cpu_data_manager_awready),                           //                    .awready
		.data_manager_wdata           (niosv_g_cpu_data_manager_wdata),                             //                    .wdata
		.data_manager_wstrb           (niosv_g_cpu_data_manager_wstrb),                             //                    .wstrb
		.data_manager_wlast           (niosv_g_cpu_data_manager_wlast),                             //                    .wlast
		.data_manager_wvalid          (niosv_g_cpu_data_manager_wvalid),                            //                    .wvalid
		.data_manager_wready          (niosv_g_cpu_data_manager_wready),                            //                    .wready
		.data_manager_bresp           (niosv_g_cpu_data_manager_bresp),                             //                    .bresp
		.data_manager_bvalid          (niosv_g_cpu_data_manager_bvalid),                            //                    .bvalid
		.data_manager_bready          (niosv_g_cpu_data_manager_bready),                            //                    .bready
		.data_manager_araddr          (niosv_g_cpu_data_manager_araddr),                            //                    .araddr
		.data_manager_arsize          (niosv_g_cpu_data_manager_arsize),                            //                    .arsize
		.data_manager_arlen           (niosv_g_cpu_data_manager_arlen),                             //                    .arlen
		.data_manager_arprot          (niosv_g_cpu_data_manager_arprot),                            //                    .arprot
		.data_manager_arvalid         (niosv_g_cpu_data_manager_arvalid),                           //                    .arvalid
		.data_manager_arready         (niosv_g_cpu_data_manager_arready),                           //                    .arready
		.data_manager_rdata           (niosv_g_cpu_data_manager_rdata),                             //                    .rdata
		.data_manager_rresp           (niosv_g_cpu_data_manager_rresp),                             //                    .rresp
		.data_manager_rvalid          (niosv_g_cpu_data_manager_rvalid),                            //                    .rvalid
		.data_manager_rlast           (niosv_g_cpu_data_manager_rlast),                             //                    .rlast
		.data_manager_rready          (niosv_g_cpu_data_manager_rready),                            //                    .rready
		.timer_sw_agent_write         (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_write),         //      timer_sw_agent.write
		.timer_sw_agent_writedata     (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_writedata),     //                    .writedata
		.timer_sw_agent_byteenable    (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_byteenable),    //                    .byteenable
		.timer_sw_agent_address       (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_address),       //                    .address
		.timer_sw_agent_read          (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_read),          //                    .read
		.timer_sw_agent_readdata      (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_readdata),      //                    .readdata
		.timer_sw_agent_readdatavalid (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_readdatavalid), //                    .readdatavalid
		.timer_sw_agent_waitrequest   (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_waitrequest),   //                    .waitrequest
		.dm_agent_write               (mm_interconnect_0_niosv_g_cpu_dm_agent_write),               //            dm_agent.write
		.dm_agent_writedata           (mm_interconnect_0_niosv_g_cpu_dm_agent_writedata),           //                    .writedata
		.dm_agent_address             (mm_interconnect_0_niosv_g_cpu_dm_agent_address),             //                    .address
		.dm_agent_read                (mm_interconnect_0_niosv_g_cpu_dm_agent_read),                //                    .read
		.dm_agent_readdata            (mm_interconnect_0_niosv_g_cpu_dm_agent_readdata),            //                    .readdata
		.dm_agent_readdatavalid       (mm_interconnect_0_niosv_g_cpu_dm_agent_readdatavalid),       //                    .readdatavalid
		.dm_agent_waitrequest         (mm_interconnect_0_niosv_g_cpu_dm_agent_waitrequest),         //                    .waitrequest
		.instruction_tcs1_awaddr      (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awaddr),      //    instruction_tcs1.awaddr
		.instruction_tcs1_awprot      (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awprot),      //                    .awprot
		.instruction_tcs1_awvalid     (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awvalid),     //                    .awvalid
		.instruction_tcs1_awready     (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awready),     //                    .awready
		.instruction_tcs1_wdata       (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wdata),       //                    .wdata
		.instruction_tcs1_wstrb       (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wstrb),       //                    .wstrb
		.instruction_tcs1_wvalid      (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wvalid),      //                    .wvalid
		.instruction_tcs1_wready      (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wready),      //                    .wready
		.instruction_tcs1_bresp       (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_bresp),       //                    .bresp
		.instruction_tcs1_bvalid      (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_bvalid),      //                    .bvalid
		.instruction_tcs1_bready      (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_bready),      //                    .bready
		.instruction_tcs1_araddr      (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_araddr),      //                    .araddr
		.instruction_tcs1_arprot      (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_arprot),      //                    .arprot
		.instruction_tcs1_arvalid     (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_arvalid),     //                    .arvalid
		.instruction_tcs1_arready     (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_arready),     //                    .arready
		.instruction_tcs1_rdata       (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rdata),       //                    .rdata
		.instruction_tcs1_rresp       (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rresp),       //                    .rresp
		.instruction_tcs1_rvalid      (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rvalid),      //                    .rvalid
		.instruction_tcs1_rready      (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rready),      //                    .rready
		.data_tcs1_awaddr             (mm_interconnect_0_niosv_g_cpu_data_tcs1_awaddr),             //           data_tcs1.awaddr
		.data_tcs1_awprot             (mm_interconnect_0_niosv_g_cpu_data_tcs1_awprot),             //                    .awprot
		.data_tcs1_awvalid            (mm_interconnect_0_niosv_g_cpu_data_tcs1_awvalid),            //                    .awvalid
		.data_tcs1_awready            (mm_interconnect_0_niosv_g_cpu_data_tcs1_awready),            //                    .awready
		.data_tcs1_wdata              (mm_interconnect_0_niosv_g_cpu_data_tcs1_wdata),              //                    .wdata
		.data_tcs1_wstrb              (mm_interconnect_0_niosv_g_cpu_data_tcs1_wstrb),              //                    .wstrb
		.data_tcs1_wvalid             (mm_interconnect_0_niosv_g_cpu_data_tcs1_wvalid),             //                    .wvalid
		.data_tcs1_wready             (mm_interconnect_0_niosv_g_cpu_data_tcs1_wready),             //                    .wready
		.data_tcs1_bresp              (mm_interconnect_0_niosv_g_cpu_data_tcs1_bresp),              //                    .bresp
		.data_tcs1_bvalid             (mm_interconnect_0_niosv_g_cpu_data_tcs1_bvalid),             //                    .bvalid
		.data_tcs1_bready             (mm_interconnect_0_niosv_g_cpu_data_tcs1_bready),             //                    .bready
		.data_tcs1_araddr             (mm_interconnect_0_niosv_g_cpu_data_tcs1_araddr),             //                    .araddr
		.data_tcs1_arprot             (mm_interconnect_0_niosv_g_cpu_data_tcs1_arprot),             //                    .arprot
		.data_tcs1_arvalid            (mm_interconnect_0_niosv_g_cpu_data_tcs1_arvalid),            //                    .arvalid
		.data_tcs1_arready            (mm_interconnect_0_niosv_g_cpu_data_tcs1_arready),            //                    .arready
		.data_tcs1_rdata              (mm_interconnect_0_niosv_g_cpu_data_tcs1_rdata),              //                    .rdata
		.data_tcs1_rresp              (mm_interconnect_0_niosv_g_cpu_data_tcs1_rresp),              //                    .rresp
		.data_tcs1_rvalid             (mm_interconnect_0_niosv_g_cpu_data_tcs1_rvalid),             //                    .rvalid
		.data_tcs1_rready             (mm_interconnect_0_niosv_g_cpu_data_tcs1_rready)              //                    .rready
	);

	NIOSV_G_SOC_SERIAL_UART_COM serial_uart_com (
		.clk           (altpll_clks_c0_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                //               reset.reset_n
		.address       (mm_interconnect_0_serial_uart_com_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_serial_uart_com_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_serial_uart_com_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_serial_uart_com_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_serial_uart_com_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_serial_uart_com_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_serial_uart_com_s1_readdata),      //                    .readdata
		.rxd           (serial_uart_com_externals_rxd),                      // external_connection.export
		.txd           (serial_uart_com_externals_txd),                      //                    .export
		.irq           (irq_mapper_receiver2_irq)                            //                 irq.irq
	);

	NIOSV_G_SOC_SOC_SYS_ID soc_sys_id (
		.clock    (altpll_clks_c0_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_soc_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_soc_sys_id_control_slave_address)   //              .address
	);

	NIOSV_G_SOC_mm_interconnect_0 mm_interconnect_0 (
		.NIOSV_G_CPU_data_manager_awaddr                               (niosv_g_cpu_data_manager_awaddr),                                    //                                NIOSV_G_CPU_data_manager.awaddr
		.NIOSV_G_CPU_data_manager_awlen                                (niosv_g_cpu_data_manager_awlen),                                     //                                                        .awlen
		.NIOSV_G_CPU_data_manager_awsize                               (niosv_g_cpu_data_manager_awsize),                                    //                                                        .awsize
		.NIOSV_G_CPU_data_manager_awprot                               (niosv_g_cpu_data_manager_awprot),                                    //                                                        .awprot
		.NIOSV_G_CPU_data_manager_awvalid                              (niosv_g_cpu_data_manager_awvalid),                                   //                                                        .awvalid
		.NIOSV_G_CPU_data_manager_awready                              (niosv_g_cpu_data_manager_awready),                                   //                                                        .awready
		.NIOSV_G_CPU_data_manager_wdata                                (niosv_g_cpu_data_manager_wdata),                                     //                                                        .wdata
		.NIOSV_G_CPU_data_manager_wstrb                                (niosv_g_cpu_data_manager_wstrb),                                     //                                                        .wstrb
		.NIOSV_G_CPU_data_manager_wlast                                (niosv_g_cpu_data_manager_wlast),                                     //                                                        .wlast
		.NIOSV_G_CPU_data_manager_wvalid                               (niosv_g_cpu_data_manager_wvalid),                                    //                                                        .wvalid
		.NIOSV_G_CPU_data_manager_wready                               (niosv_g_cpu_data_manager_wready),                                    //                                                        .wready
		.NIOSV_G_CPU_data_manager_bresp                                (niosv_g_cpu_data_manager_bresp),                                     //                                                        .bresp
		.NIOSV_G_CPU_data_manager_bvalid                               (niosv_g_cpu_data_manager_bvalid),                                    //                                                        .bvalid
		.NIOSV_G_CPU_data_manager_bready                               (niosv_g_cpu_data_manager_bready),                                    //                                                        .bready
		.NIOSV_G_CPU_data_manager_araddr                               (niosv_g_cpu_data_manager_araddr),                                    //                                                        .araddr
		.NIOSV_G_CPU_data_manager_arlen                                (niosv_g_cpu_data_manager_arlen),                                     //                                                        .arlen
		.NIOSV_G_CPU_data_manager_arsize                               (niosv_g_cpu_data_manager_arsize),                                    //                                                        .arsize
		.NIOSV_G_CPU_data_manager_arprot                               (niosv_g_cpu_data_manager_arprot),                                    //                                                        .arprot
		.NIOSV_G_CPU_data_manager_arvalid                              (niosv_g_cpu_data_manager_arvalid),                                   //                                                        .arvalid
		.NIOSV_G_CPU_data_manager_arready                              (niosv_g_cpu_data_manager_arready),                                   //                                                        .arready
		.NIOSV_G_CPU_data_manager_rdata                                (niosv_g_cpu_data_manager_rdata),                                     //                                                        .rdata
		.NIOSV_G_CPU_data_manager_rresp                                (niosv_g_cpu_data_manager_rresp),                                     //                                                        .rresp
		.NIOSV_G_CPU_data_manager_rlast                                (niosv_g_cpu_data_manager_rlast),                                     //                                                        .rlast
		.NIOSV_G_CPU_data_manager_rvalid                               (niosv_g_cpu_data_manager_rvalid),                                    //                                                        .rvalid
		.NIOSV_G_CPU_data_manager_rready                               (niosv_g_cpu_data_manager_rready),                                    //                                                        .rready
		.NIOSV_G_CPU_data_tcs1_awaddr                                  (mm_interconnect_0_niosv_g_cpu_data_tcs1_awaddr),                     //                                   NIOSV_G_CPU_data_tcs1.awaddr
		.NIOSV_G_CPU_data_tcs1_awprot                                  (mm_interconnect_0_niosv_g_cpu_data_tcs1_awprot),                     //                                                        .awprot
		.NIOSV_G_CPU_data_tcs1_awvalid                                 (mm_interconnect_0_niosv_g_cpu_data_tcs1_awvalid),                    //                                                        .awvalid
		.NIOSV_G_CPU_data_tcs1_awready                                 (mm_interconnect_0_niosv_g_cpu_data_tcs1_awready),                    //                                                        .awready
		.NIOSV_G_CPU_data_tcs1_wdata                                   (mm_interconnect_0_niosv_g_cpu_data_tcs1_wdata),                      //                                                        .wdata
		.NIOSV_G_CPU_data_tcs1_wstrb                                   (mm_interconnect_0_niosv_g_cpu_data_tcs1_wstrb),                      //                                                        .wstrb
		.NIOSV_G_CPU_data_tcs1_wvalid                                  (mm_interconnect_0_niosv_g_cpu_data_tcs1_wvalid),                     //                                                        .wvalid
		.NIOSV_G_CPU_data_tcs1_wready                                  (mm_interconnect_0_niosv_g_cpu_data_tcs1_wready),                     //                                                        .wready
		.NIOSV_G_CPU_data_tcs1_bresp                                   (mm_interconnect_0_niosv_g_cpu_data_tcs1_bresp),                      //                                                        .bresp
		.NIOSV_G_CPU_data_tcs1_bvalid                                  (mm_interconnect_0_niosv_g_cpu_data_tcs1_bvalid),                     //                                                        .bvalid
		.NIOSV_G_CPU_data_tcs1_bready                                  (mm_interconnect_0_niosv_g_cpu_data_tcs1_bready),                     //                                                        .bready
		.NIOSV_G_CPU_data_tcs1_araddr                                  (mm_interconnect_0_niosv_g_cpu_data_tcs1_araddr),                     //                                                        .araddr
		.NIOSV_G_CPU_data_tcs1_arprot                                  (mm_interconnect_0_niosv_g_cpu_data_tcs1_arprot),                     //                                                        .arprot
		.NIOSV_G_CPU_data_tcs1_arvalid                                 (mm_interconnect_0_niosv_g_cpu_data_tcs1_arvalid),                    //                                                        .arvalid
		.NIOSV_G_CPU_data_tcs1_arready                                 (mm_interconnect_0_niosv_g_cpu_data_tcs1_arready),                    //                                                        .arready
		.NIOSV_G_CPU_data_tcs1_rdata                                   (mm_interconnect_0_niosv_g_cpu_data_tcs1_rdata),                      //                                                        .rdata
		.NIOSV_G_CPU_data_tcs1_rresp                                   (mm_interconnect_0_niosv_g_cpu_data_tcs1_rresp),                      //                                                        .rresp
		.NIOSV_G_CPU_data_tcs1_rvalid                                  (mm_interconnect_0_niosv_g_cpu_data_tcs1_rvalid),                     //                                                        .rvalid
		.NIOSV_G_CPU_data_tcs1_rready                                  (mm_interconnect_0_niosv_g_cpu_data_tcs1_rready),                     //                                                        .rready
		.NIOSV_G_CPU_instruction_manager_awaddr                        (niosv_g_cpu_instruction_manager_awaddr),                             //                         NIOSV_G_CPU_instruction_manager.awaddr
		.NIOSV_G_CPU_instruction_manager_awlen                         (niosv_g_cpu_instruction_manager_awlen),                              //                                                        .awlen
		.NIOSV_G_CPU_instruction_manager_awsize                        (niosv_g_cpu_instruction_manager_awsize),                             //                                                        .awsize
		.NIOSV_G_CPU_instruction_manager_awburst                       (niosv_g_cpu_instruction_manager_awburst),                            //                                                        .awburst
		.NIOSV_G_CPU_instruction_manager_awprot                        (niosv_g_cpu_instruction_manager_awprot),                             //                                                        .awprot
		.NIOSV_G_CPU_instruction_manager_awvalid                       (niosv_g_cpu_instruction_manager_awvalid),                            //                                                        .awvalid
		.NIOSV_G_CPU_instruction_manager_awready                       (niosv_g_cpu_instruction_manager_awready),                            //                                                        .awready
		.NIOSV_G_CPU_instruction_manager_wdata                         (niosv_g_cpu_instruction_manager_wdata),                              //                                                        .wdata
		.NIOSV_G_CPU_instruction_manager_wstrb                         (niosv_g_cpu_instruction_manager_wstrb),                              //                                                        .wstrb
		.NIOSV_G_CPU_instruction_manager_wlast                         (niosv_g_cpu_instruction_manager_wlast),                              //                                                        .wlast
		.NIOSV_G_CPU_instruction_manager_wvalid                        (niosv_g_cpu_instruction_manager_wvalid),                             //                                                        .wvalid
		.NIOSV_G_CPU_instruction_manager_wready                        (niosv_g_cpu_instruction_manager_wready),                             //                                                        .wready
		.NIOSV_G_CPU_instruction_manager_bresp                         (niosv_g_cpu_instruction_manager_bresp),                              //                                                        .bresp
		.NIOSV_G_CPU_instruction_manager_bvalid                        (niosv_g_cpu_instruction_manager_bvalid),                             //                                                        .bvalid
		.NIOSV_G_CPU_instruction_manager_bready                        (niosv_g_cpu_instruction_manager_bready),                             //                                                        .bready
		.NIOSV_G_CPU_instruction_manager_araddr                        (niosv_g_cpu_instruction_manager_araddr),                             //                                                        .araddr
		.NIOSV_G_CPU_instruction_manager_arlen                         (niosv_g_cpu_instruction_manager_arlen),                              //                                                        .arlen
		.NIOSV_G_CPU_instruction_manager_arsize                        (niosv_g_cpu_instruction_manager_arsize),                             //                                                        .arsize
		.NIOSV_G_CPU_instruction_manager_arburst                       (niosv_g_cpu_instruction_manager_arburst),                            //                                                        .arburst
		.NIOSV_G_CPU_instruction_manager_arprot                        (niosv_g_cpu_instruction_manager_arprot),                             //                                                        .arprot
		.NIOSV_G_CPU_instruction_manager_arvalid                       (niosv_g_cpu_instruction_manager_arvalid),                            //                                                        .arvalid
		.NIOSV_G_CPU_instruction_manager_arready                       (niosv_g_cpu_instruction_manager_arready),                            //                                                        .arready
		.NIOSV_G_CPU_instruction_manager_rdata                         (niosv_g_cpu_instruction_manager_rdata),                              //                                                        .rdata
		.NIOSV_G_CPU_instruction_manager_rresp                         (niosv_g_cpu_instruction_manager_rresp),                              //                                                        .rresp
		.NIOSV_G_CPU_instruction_manager_rlast                         (niosv_g_cpu_instruction_manager_rlast),                              //                                                        .rlast
		.NIOSV_G_CPU_instruction_manager_rvalid                        (niosv_g_cpu_instruction_manager_rvalid),                             //                                                        .rvalid
		.NIOSV_G_CPU_instruction_manager_rready                        (niosv_g_cpu_instruction_manager_rready),                             //                                                        .rready
		.NIOSV_G_CPU_instruction_tcs1_awaddr                           (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awaddr),              //                            NIOSV_G_CPU_instruction_tcs1.awaddr
		.NIOSV_G_CPU_instruction_tcs1_awprot                           (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awprot),              //                                                        .awprot
		.NIOSV_G_CPU_instruction_tcs1_awvalid                          (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awvalid),             //                                                        .awvalid
		.NIOSV_G_CPU_instruction_tcs1_awready                          (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_awready),             //                                                        .awready
		.NIOSV_G_CPU_instruction_tcs1_wdata                            (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wdata),               //                                                        .wdata
		.NIOSV_G_CPU_instruction_tcs1_wstrb                            (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wstrb),               //                                                        .wstrb
		.NIOSV_G_CPU_instruction_tcs1_wvalid                           (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wvalid),              //                                                        .wvalid
		.NIOSV_G_CPU_instruction_tcs1_wready                           (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_wready),              //                                                        .wready
		.NIOSV_G_CPU_instruction_tcs1_bresp                            (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_bresp),               //                                                        .bresp
		.NIOSV_G_CPU_instruction_tcs1_bvalid                           (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_bvalid),              //                                                        .bvalid
		.NIOSV_G_CPU_instruction_tcs1_bready                           (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_bready),              //                                                        .bready
		.NIOSV_G_CPU_instruction_tcs1_araddr                           (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_araddr),              //                                                        .araddr
		.NIOSV_G_CPU_instruction_tcs1_arprot                           (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_arprot),              //                                                        .arprot
		.NIOSV_G_CPU_instruction_tcs1_arvalid                          (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_arvalid),             //                                                        .arvalid
		.NIOSV_G_CPU_instruction_tcs1_arready                          (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_arready),             //                                                        .arready
		.NIOSV_G_CPU_instruction_tcs1_rdata                            (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rdata),               //                                                        .rdata
		.NIOSV_G_CPU_instruction_tcs1_rresp                            (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rresp),               //                                                        .rresp
		.NIOSV_G_CPU_instruction_tcs1_rvalid                           (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rvalid),              //                                                        .rvalid
		.NIOSV_G_CPU_instruction_tcs1_rready                           (mm_interconnect_0_niosv_g_cpu_instruction_tcs1_rready),              //                                                        .rready
		.ALTPLL_CLKS_c0_clk                                            (altpll_clks_c0_clk),                                                 //                                          ALTPLL_CLKS_c0.clk
		.ALTPLL_CLKS_c2_clk                                            (altpll_clks_c2_clk),                                                 //                                          ALTPLL_CLKS_c2.clk
		.CLOCK_BRIDGE_IN_out_clk_clk                                   (clock_bridge_in_clk_clk),                                            //                                 CLOCK_BRIDGE_IN_out_clk.clk
		.ALTPLL_CLKS_inclk_interface_reset_reset_bridge_in_reset_reset (~reset_bridge_in_reset_n_reset_n),                                   // ALTPLL_CLKS_inclk_interface_reset_reset_bridge_in_reset.reset
		.EPCS_FLASH_CONTROLLER_PROG_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                                     //  EPCS_FLASH_CONTROLLER_PROG_reset_reset_bridge_in_reset.reset
		.NIOSV_G_CPU_reset_reset_bridge_in_reset_reset                 (rst_controller_001_reset_out_reset),                                 //                 NIOSV_G_CPU_reset_reset_bridge_in_reset.reset
		.ALTPLL_CLKS_pll_slave_address                                 (mm_interconnect_0_altpll_clks_pll_slave_address),                    //                                   ALTPLL_CLKS_pll_slave.address
		.ALTPLL_CLKS_pll_slave_write                                   (mm_interconnect_0_altpll_clks_pll_slave_write),                      //                                                        .write
		.ALTPLL_CLKS_pll_slave_read                                    (mm_interconnect_0_altpll_clks_pll_slave_read),                       //                                                        .read
		.ALTPLL_CLKS_pll_slave_readdata                                (mm_interconnect_0_altpll_clks_pll_slave_readdata),                   //                                                        .readdata
		.ALTPLL_CLKS_pll_slave_writedata                               (mm_interconnect_0_altpll_clks_pll_slave_writedata),                  //                                                        .writedata
		.EPCS_FLASH_CONTROLLER_PROG_avl_csr_address                    (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_address),       //                      EPCS_FLASH_CONTROLLER_PROG_avl_csr.address
		.EPCS_FLASH_CONTROLLER_PROG_avl_csr_write                      (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_write),         //                                                        .write
		.EPCS_FLASH_CONTROLLER_PROG_avl_csr_read                       (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_read),          //                                                        .read
		.EPCS_FLASH_CONTROLLER_PROG_avl_csr_readdata                   (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_readdata),      //                                                        .readdata
		.EPCS_FLASH_CONTROLLER_PROG_avl_csr_writedata                  (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_writedata),     //                                                        .writedata
		.EPCS_FLASH_CONTROLLER_PROG_avl_csr_readdatavalid              (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_readdatavalid), //                                                        .readdatavalid
		.EPCS_FLASH_CONTROLLER_PROG_avl_csr_waitrequest                (mm_interconnect_0_epcs_flash_controller_prog_avl_csr_waitrequest),   //                                                        .waitrequest
		.EPCS_FLASH_CONTROLLER_PROG_avl_mem_address                    (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_address),       //                      EPCS_FLASH_CONTROLLER_PROG_avl_mem.address
		.EPCS_FLASH_CONTROLLER_PROG_avl_mem_write                      (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_write),         //                                                        .write
		.EPCS_FLASH_CONTROLLER_PROG_avl_mem_read                       (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_read),          //                                                        .read
		.EPCS_FLASH_CONTROLLER_PROG_avl_mem_readdata                   (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_readdata),      //                                                        .readdata
		.EPCS_FLASH_CONTROLLER_PROG_avl_mem_writedata                  (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_writedata),     //                                                        .writedata
		.EPCS_FLASH_CONTROLLER_PROG_avl_mem_burstcount                 (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_burstcount),    //                                                        .burstcount
		.EPCS_FLASH_CONTROLLER_PROG_avl_mem_byteenable                 (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_byteenable),    //                                                        .byteenable
		.EPCS_FLASH_CONTROLLER_PROG_avl_mem_readdatavalid              (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_readdatavalid), //                                                        .readdatavalid
		.EPCS_FLASH_CONTROLLER_PROG_avl_mem_waitrequest                (mm_interconnect_0_epcs_flash_controller_prog_avl_mem_waitrequest),   //                                                        .waitrequest
		.GPI0_BTN_s1_address                                           (mm_interconnect_0_gpi0_btn_s1_address),                              //                                             GPI0_BTN_s1.address
		.GPI0_BTN_s1_write                                             (mm_interconnect_0_gpi0_btn_s1_write),                                //                                                        .write
		.GPI0_BTN_s1_readdata                                          (mm_interconnect_0_gpi0_btn_s1_readdata),                             //                                                        .readdata
		.GPI0_BTN_s1_writedata                                         (mm_interconnect_0_gpi0_btn_s1_writedata),                            //                                                        .writedata
		.GPI0_BTN_s1_chipselect                                        (mm_interconnect_0_gpi0_btn_s1_chipselect),                           //                                                        .chipselect
		.GPI1_DIPSW_s1_address                                         (mm_interconnect_0_gpi1_dipsw_s1_address),                            //                                           GPI1_DIPSW_s1.address
		.GPI1_DIPSW_s1_write                                           (mm_interconnect_0_gpi1_dipsw_s1_write),                              //                                                        .write
		.GPI1_DIPSW_s1_readdata                                        (mm_interconnect_0_gpi1_dipsw_s1_readdata),                           //                                                        .readdata
		.GPI1_DIPSW_s1_writedata                                       (mm_interconnect_0_gpi1_dipsw_s1_writedata),                          //                                                        .writedata
		.GPI1_DIPSW_s1_chipselect                                      (mm_interconnect_0_gpi1_dipsw_s1_chipselect),                         //                                                        .chipselect
		.GPO2_LEDG_s1_address                                          (mm_interconnect_0_gpo2_ledg_s1_address),                             //                                            GPO2_LEDG_s1.address
		.GPO2_LEDG_s1_write                                            (mm_interconnect_0_gpo2_ledg_s1_write),                               //                                                        .write
		.GPO2_LEDG_s1_readdata                                         (mm_interconnect_0_gpo2_ledg_s1_readdata),                            //                                                        .readdata
		.GPO2_LEDG_s1_writedata                                        (mm_interconnect_0_gpo2_ledg_s1_writedata),                           //                                                        .writedata
		.GPO2_LEDG_s1_chipselect                                       (mm_interconnect_0_gpo2_ledg_s1_chipselect),                          //                                                        .chipselect
		.JTAG_UART_COM_avalon_jtag_slave_address                       (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_address),          //                         JTAG_UART_COM_avalon_jtag_slave.address
		.JTAG_UART_COM_avalon_jtag_slave_write                         (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_write),            //                                                        .write
		.JTAG_UART_COM_avalon_jtag_slave_read                          (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_read),             //                                                        .read
		.JTAG_UART_COM_avalon_jtag_slave_readdata                      (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_readdata),         //                                                        .readdata
		.JTAG_UART_COM_avalon_jtag_slave_writedata                     (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_writedata),        //                                                        .writedata
		.JTAG_UART_COM_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_waitrequest),      //                                                        .waitrequest
		.JTAG_UART_COM_avalon_jtag_slave_chipselect                    (mm_interconnect_0_jtag_uart_com_avalon_jtag_slave_chipselect),       //                                                        .chipselect
		.NIOSV_G_CPU_dm_agent_address                                  (mm_interconnect_0_niosv_g_cpu_dm_agent_address),                     //                                    NIOSV_G_CPU_dm_agent.address
		.NIOSV_G_CPU_dm_agent_write                                    (mm_interconnect_0_niosv_g_cpu_dm_agent_write),                       //                                                        .write
		.NIOSV_G_CPU_dm_agent_read                                     (mm_interconnect_0_niosv_g_cpu_dm_agent_read),                        //                                                        .read
		.NIOSV_G_CPU_dm_agent_readdata                                 (mm_interconnect_0_niosv_g_cpu_dm_agent_readdata),                    //                                                        .readdata
		.NIOSV_G_CPU_dm_agent_writedata                                (mm_interconnect_0_niosv_g_cpu_dm_agent_writedata),                   //                                                        .writedata
		.NIOSV_G_CPU_dm_agent_readdatavalid                            (mm_interconnect_0_niosv_g_cpu_dm_agent_readdatavalid),               //                                                        .readdatavalid
		.NIOSV_G_CPU_dm_agent_waitrequest                              (mm_interconnect_0_niosv_g_cpu_dm_agent_waitrequest),                 //                                                        .waitrequest
		.NIOSV_G_CPU_timer_sw_agent_address                            (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_address),               //                              NIOSV_G_CPU_timer_sw_agent.address
		.NIOSV_G_CPU_timer_sw_agent_write                              (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_write),                 //                                                        .write
		.NIOSV_G_CPU_timer_sw_agent_read                               (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_read),                  //                                                        .read
		.NIOSV_G_CPU_timer_sw_agent_readdata                           (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_readdata),              //                                                        .readdata
		.NIOSV_G_CPU_timer_sw_agent_writedata                          (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_writedata),             //                                                        .writedata
		.NIOSV_G_CPU_timer_sw_agent_byteenable                         (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_byteenable),            //                                                        .byteenable
		.NIOSV_G_CPU_timer_sw_agent_readdatavalid                      (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_readdatavalid),         //                                                        .readdatavalid
		.NIOSV_G_CPU_timer_sw_agent_waitrequest                        (mm_interconnect_0_niosv_g_cpu_timer_sw_agent_waitrequest),           //                                                        .waitrequest
		.SERIAL_UART_COM_s1_address                                    (mm_interconnect_0_serial_uart_com_s1_address),                       //                                      SERIAL_UART_COM_s1.address
		.SERIAL_UART_COM_s1_write                                      (mm_interconnect_0_serial_uart_com_s1_write),                         //                                                        .write
		.SERIAL_UART_COM_s1_read                                       (mm_interconnect_0_serial_uart_com_s1_read),                          //                                                        .read
		.SERIAL_UART_COM_s1_readdata                                   (mm_interconnect_0_serial_uart_com_s1_readdata),                      //                                                        .readdata
		.SERIAL_UART_COM_s1_writedata                                  (mm_interconnect_0_serial_uart_com_s1_writedata),                     //                                                        .writedata
		.SERIAL_UART_COM_s1_begintransfer                              (mm_interconnect_0_serial_uart_com_s1_begintransfer),                 //                                                        .begintransfer
		.SERIAL_UART_COM_s1_chipselect                                 (mm_interconnect_0_serial_uart_com_s1_chipselect),                    //                                                        .chipselect
		.SOC_SYS_ID_control_slave_address                              (mm_interconnect_0_soc_sys_id_control_slave_address),                 //                                SOC_SYS_ID_control_slave.address
		.SOC_SYS_ID_control_slave_readdata                             (mm_interconnect_0_soc_sys_id_control_slave_readdata)                 //                                                        .readdata
	);

	NIOSV_G_SOC_irq_mapper irq_mapper (
		.clk           (altpll_clks_c0_clk),                 //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (niosv_g_cpu_platform_irq_rx_irq)     //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_clks_c2_clk),                 //       receiver_clk.clk
		.sender_clk     (altpll_clks_c0_clk),                 //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_bridge_in_reset_n_reset_n), // reset_in0.reset
		.clk            (altpll_clks_c2_clk),               //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                 // (terminated)
		.reset_req_in0  (1'b0),                             // (terminated)
		.reset_in1      (1'b0),                             // (terminated)
		.reset_req_in1  (1'b0),                             // (terminated)
		.reset_in2      (1'b0),                             // (terminated)
		.reset_req_in2  (1'b0),                             // (terminated)
		.reset_in3      (1'b0),                             // (terminated)
		.reset_req_in3  (1'b0),                             // (terminated)
		.reset_in4      (1'b0),                             // (terminated)
		.reset_req_in4  (1'b0),                             // (terminated)
		.reset_in5      (1'b0),                             // (terminated)
		.reset_req_in5  (1'b0),                             // (terminated)
		.reset_in6      (1'b0),                             // (terminated)
		.reset_req_in6  (1'b0),                             // (terminated)
		.reset_in7      (1'b0),                             // (terminated)
		.reset_req_in7  (1'b0),                             // (terminated)
		.reset_in8      (1'b0),                             // (terminated)
		.reset_req_in8  (1'b0),                             // (terminated)
		.reset_in9      (1'b0),                             // (terminated)
		.reset_req_in9  (1'b0),                             // (terminated)
		.reset_in10     (1'b0),                             // (terminated)
		.reset_req_in10 (1'b0),                             // (terminated)
		.reset_in11     (1'b0),                             // (terminated)
		.reset_req_in11 (1'b0),                             // (terminated)
		.reset_in12     (1'b0),                             // (terminated)
		.reset_req_in12 (1'b0),                             // (terminated)
		.reset_in13     (1'b0),                             // (terminated)
		.reset_req_in13 (1'b0),                             // (terminated)
		.reset_in14     (1'b0),                             // (terminated)
		.reset_req_in14 (1'b0),                             // (terminated)
		.reset_in15     (1'b0),                             // (terminated)
		.reset_req_in15 (1'b0)                              // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_bridge_in_reset_n_reset_n),   // reset_in0.reset
		.clk            (altpll_clks_c0_clk),                 //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
