��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a�����{������#��j��{��	?+�g��-��"XSʌb������;�b���/��.v���9�Cr� x�B ��q���mL)�-�"6|��hHwg��	��j������猽?�����?�__��n$ԗ�����NÀ�-
�R�6�d��v�����t;��df�!�+#G��Բ��87E�1�R�x��)O�+�w�v\�A�B�i�y_7V)�5`�@uș����J��E��9zuS�H5U���	�#�%����BV��95[� Y����J�g�qfKD<������ �_.?�ǉE��1�?�1+��P|�-�D����4��Kt~v�v-�k��%i^ո�Z;�Ƥ�������̭�^
;'�}6Y��#e����5������M�;v�	�m����v�UB��� ���tj�
��p��e�#��FrSŶ�3�,nu�y����뻬��(V^1Zv��6�W��~tb��Pz�SV�N��.R�ܕl~�Uq/�]���+ɫs�d�'��}F�Yh���t70�.$��hŏ���t��<ޙ�*����1��Ta�E������ ϶|���9��NF	\�B�A�n�{\���J��ˬ�fW����Br��{%����q���@F#�*��ә�֥\�[$)T�kn?Ї����v�d23�E��8'D�Q��6h*�Iq7�!��c��;�MklK��=6^s;�v��¢���[���'�V��1�wXD���!W��{什xeq����Ȓ�~#�v	�����P%��B���x��_��x���R�^����x9��UD��#��U����o4t7~�p��)��}B*>X�Иɋa��\�c�TãB�������ڻUG;�a��H��)2�������A& ���j�dSI���̀J�,�m6�y%�S̹*	c�$׍��dy��S�2v�?i�mK��y.F�_+	��g,5� ��2�ɖ�#��H8yi�G�;�w'Ҷ�C]Z�$�)Ä+�t	.:������!���2�L[��A�υj��/�+��y�-���@Y+С��}�Q|D�(C س�G^���
]��0&룖)����6�v���LP�ըdxic� 
�zR
�w�3��������|��ꍝd��h)�k��\����^s9ubl�Sw�Qы��j���+�MC)����W�A/g�Z���d���N��ԑ��q�;����G�_�0��EJ�{X�l2n����L�r����!�"���B$O�Z���{����)���y�ML�P��QH�N�q�&�9:
a)���$���|����`٘��%���q��X0G�o����%���Q��~E�דXMeq+��1�u2ҪP`o�7tY�z�%'�@�(_=I	^��FkB�>��0L��IR�����u�G��@!7�ԷA9�N�}��c��l�-�9��P��^o !�Q[E��I8�����?�$_�RI���^�R̶@}�2< |��_���T]��S�=t$ux/� lX����|.� �2���2��?o��hW�-�"p���Eo0O��aV"��	�s� "U_c�$��XqiX�B)�eF���+4�?�+iUg���Ӳf��,f�S��}瑏V�?z�R���X��Q�g�<2z3
ٞxl�Ƣ���q���/LH<b�oP��50��1��ӧmg��D����{�W�@_Z	��pDq�"�A�O��������̅2B��7mr&�U�&rD��ˡ�P�
j|�^�10����\�r YR���ꬺl���	r�,�Ge�y�gHd��J�Jn�ߘ���,z�n��x��ߓ�n�a�T�S�}k��x����MG�L�:��y�Pl��B���V���y��vMkwF��G܆G^�2%��"��18[J�ƌ�:��5��Q��S(��kׄf8EYX�� @
�2���kb��.��]��[�_��
ǶW�D�g,�"��ۓ�3~YSvFb�4ikc���r��w=�$3qD���Ґ�?No��>�
0祾_�OMK.�/4n{~�~G�������T�G*8�%�j�W��3w�w8�Aʫ�^0��{N��0 (�>~5�=f%E����#�f��z��`�H���b���V�:'R�͝�u�5����G�d���P���H՞o	���8k�-��>�ӌ<����<sd�)gr��/ ���z�Vע*YB�!�C�RR��@�ys��\�Ag��O�oo��u�ҹC�"�#�!�/�U���!vm*�����4X��8݋c��{81��rJ�;��C�쭤�!A��{+�h���-y]k��3�Ц�?�5��Ϣ\_l]����_�_��`xז��,5���pM�F���O��G"g]�u�HR�!�Y/Չ�5���
��ƻm��"�QG�kdoLBo��'�P|÷C�2Ȧ�#D�P�J��)�ʆ���'�'���+�r���Uf_wt��X�i�M6T��"&��vI�=�,�]F�q'����.!
A�ݙz���Ѧ�7��A��?�]��Ϊ|~��n$ؔc�/7�[�b8�v@n���h0��sW���26a�������YM��M��:��Ns3}�G6� ;/0��DH�E�w�Q� S�c�W>x�r�~nN��?��#sz�Y��b��3�c㲍����;�($N�	_��&נ[�Fҫ��Y6��ٽZ�r�g]�Ww����%X$DW��q�`��xwB���j�yd����x0'�P�܎��ͧ�0�����$�ڧFΣ,8<~U��ḧ�1R}J�P7C����<(u���ܓlOd���'.c�� u�־t���MͲg�}���6`Pұ[����. []�+7sY^�8�d?a�5��3<�ú��?)+��ׄ�jI ���h *b	tY��(
�<�����/�;A,��)N�E���Ņ��%�'Qm[j]�xֽ�O��2�Ծc߼�}�����Ȁ!���-2��g���&ܒ*������@�Z����,Qց>�
R�<H4�G��:9�a�e�>i����ș!.0�j�au����.�U ���3���s5wh��-�s"Zk�,�eێ���[l�����k�����t��_L����'���l�Te�};�]�b`��O=%�x5�9a(��y��"�N6	�D� Q�rć0����pO�����j�uzo�@���ȵ�۳OQ��{��L��Fr�M �^�@�z����/@���4Ӎ@b��*3C���3�a9p��I߀�G>B���Tv�{��1��ǫG%q��q�p�a��dBj��0ď�U)��0ΎK|qz��=r�"`������������n���.���W�Ӭ�J������G�.Nqٱx���'����iv-~p���/�3�*{eK;!DA�����EM�KBʲ ���6���=?�Oy���Ħ�d��V���
],�I��]�gC�ڿ���\U���}����z} �qb�T ´*;�iJR�ޟt	�9���U`�l�_�=/��>����6{{>5	�4	�o����a�lz�[I0�k�|�,�<lr�T ���Z�������7O_�f�LO��9���i�#mF�L�4_t�ږ,�j�]��`[yɛ���C�0�s������� �R��k�CQ*~ƣs� �~<^��۴�Ӏ-���,�M�)خ��m�5����/k*�>�<�r�i������b���AG�681]�kdY��8�"��y�����"}��4�X]�����x�F�g�Jڒ1�{ւ�v�
�Z�2�:K*HUI"������z�&�a�o�:{���eJ/Ҍ�ٮ�nP�xҘ >Дd�d7edO�����@߄9dS�FT�:��M�#{���"��炋�6hTn��a�A�E�ۗ����Cv�~�x	�4��Ͼ2E�d�������&:�X)��Kscp�1���ꐡ֝hS��c3A}�B�`i*�O��>թ��!@pʴ�	�΅�3Cs��P���'׍Y���h!�{�j�P�H�/�k�QUMm�9����1�6����3���o��Wb��I8�uU���)$��Ei2֭�U��D����7|;���-/�5��r��x�����}���|,E�x�R|����g�fxu`�շ���Co|\�X4pr?���G_��ňT;:��;b9Y93��*����bi�@�����/:Ɗ#��$!�������f�8�_z���Ūi���Wj�W���?�y�k���LY�I�c���1�J�Z�H��O���)���k�Nu��,����h��z7��ζ`<�'�ä5&"�:��D+�˟!��z�+�,j���c���ؑ[$�&�'��sWG�qj�JHA�I·Yȋ������ā�x�J�U݁ؕe8��%>ǪqV��S�"*^ Lp��[�"�#��ƚL�t,�U��гK�X�=���x
䆽ga&��U�}�4�V'�x<��)�@�:/M8lÒ@,�53�dK�@�S#��v�_�>�FG!�>P��cЛQ�x���+~^�\�r0L����ÜsM�x�|;!��r>����Q�$c�T}5��_U��FT���z�f_��M��X�(5��J݆������~�� Ռ�R��0�l�\)���|�0�]���n���C&Ү�Zb-P̶G��:�/s}��h���4ߺ�جT��>X��jLp��A&���.V�VS�3�����4����l�A5{5 Ej�q�<���8��+�1��Q;�Po5Ҏ��g:�#zb��΄*�:eTC��閟�%�JC���`}ȤAEYϳs�fa�#���Ŝ��5�>�'ѱ����+�⎐GW9� �X��~%��a���M�=��xk%���c�~�)+���fb�6�+5�{L����d���_�kQ��w��~�:
πZќifk.��߄V��Kf��n5>��|�Y�Kus��R���p ��&�����"ڰ�\K;���F���j�3be���~��|�ς��6)��l;��ǯm|�P�GmS_Qb���4	)u����}$+E��F����?݃:�� q�q�?@�����L��9};�cI�@�D�~5����>�&�8��/5�hnTΩN;c4���X���R�S���T�uJgLUJ��fV�{��4�H.�(�Ї�k�Xl=!��<w\�K�`U���,�b$���O������*�@c��`�;��a��D���/����(���z�zpn�YT�z��^q�D���ok��!���O�q�Ԭ�?F��#~d�DixǶ��{�č
Ja���z� ;%2�k�{�)��ɟ�QLi����t/mE9c�ir9(���)�����s��N����TH��:c!�Ds����h���Ɉ��ځtB4�Uw(-.仡�px$��Ű��m�y�6��G��4e�Fh��6��rSo:���M����R���ZXۀϼ[NA7�����m��/�����	�M�}�b&��sq�����w�ڥC��GԱj�F�&��
ٍ�meX �N�e��4�j����y\��ۆ6Y@�9�,^ga�}�Qd�O�����0�*�
���3�����{L�j�le�'N8���ϳ�C���}R嬻��7Ę�G+�\Z����^�{��ǖAJ�p�A�E[���=�2rO��[��/[G˱>���Hs�TB��νn ��hurp��pr�Xx�q	��hDl�T���6���*�o=�mhke��Xɩ��q�n]c�P���а�_t�(^�.`�$d�t�I,s�N��/y�+DΫY���Ex��(�}3o�]!���D,||�&���˰i��r3ʔ�)�	V!bݡ��JԶmpvn����NJK����AA6tz"�V x�9��6Μ�r�����8�L�];��u�1:����Ӥ��oO��(从�@�{�g�lb��1m�
W0��Lw��ǈ���RQ�=�a�o��y�P�M�D��D�<|×m�0�*��x�_]�s����Y!���d�R7���Q5�Nh�9�}�3d�&�kJ�QLz����[7ɿ�����O��+��M�<���eqM@6YD����Ԏ��}:G�
,�ȇy��"��~H�ɹ��	9id3�x +���,߁@�9���+g��'KnA�;���(P���vih���l̇k��6tꈽ��	�����rFf��������GG��r��h��"�4ba=����?����/�FL�9�y������Wz�O�2P��B)�)`�c_�z�^3+�xq�c��5�+aU��n�[$P�a��#o�W���RP?�m��T�����bi�EW&��D �&Ɖ��c
.�Ej�7�R��R&6�����k)d~ʴ��r�}��lX 36�1�rz�n���]��p��
�N|���'�N	*����þ���Zh�]��A�}!�S��9�Yl��q<�� í�S2E�.�¸��6j��/��A@�rssWį*�V=s��CRёPp�������K�;0�*�@�?�������_*�F��_qZ
 �y���@��=U$'�O>��H#��AB~@�8u(��E6 �s�2�䴥>���RɃ������|dHoL��b,'�s���,�9s�s�s����\�ϗ����;e!4�?�/ e��V��[���X�Y�{w��Y~z�|�(��{����"��f{�}�wm��&�����mq������tV�(8���ŪU�/�Q��h�&���90MM��yd�&f��{v�����:2�IȂ"��H��[�}���fXMŐ8.�tCq��p��&����jK��itՃ+6�4Ll$7� #+�70��ȩz�0�e�Y)�@꿟frï�F��`���l��F�e)y._�Oڊ��W�E�Y��_����n��&���!�9��D5zf�=L685���"��ta=�7�i�ĵ��n3�m�~ہ��i�����T�aב���t���o4 �aҙ��P��:��0��q-�6���e�����tr�Ѳ5��R&�}INAH��Er���7�&jl����ýC�;�01�����枋g��� j���!95��L���"��2-��q\b�Y51��=k�y���S�c���uj��mu�;�.�Q�Z[��J�������wӊ�+��H��%I���H���� ��[�T6�M��q�X " �&�[������zo��!���:�aR�)�ڐ�>'!�8�����|���,���$i���y�9������6�$�f�ϯ����̖|�ޭ�At�ꕚ����h��?�H0�`�Y�u��ސ������>�$��`H�t�Г��U�~���>p@R���x�O;�s�W",��O��*�X�)���r���a�q����%ג�4�f�	z��G�~��]���%�m�j��c)�X$�m����a�	��"�7��Ƴ�_�
��m��7��3�4��w!�����i����e*��V�w�tC����D����}���9�ƌ.��Q��3\�vI��Y�hҦ*���
�KL��gQg� �Q�����
/�e�EXBY���MCts��gv�:9gn�(u�.�pP�6�`	`�_�D�������w������wZ�<��Dk	��<Q�/��~��>���QErS�2%1�.��8|��h��։IeiIM}l �l8= H���Mw�9�nP�
mz�*-�����
�3GZ2FQ �]F2�8�05��=1�jc��kC���MyQ/��	L�JT�z��%�`���Fï�+Z�z�#5�#� ��mQ{�k �>\AqB����M�+J��2͹gOʛ���H��L}�cH��x�wH̺c��[/�`�/�H�j{�7hd'��9e6G��=�s�kn��%1�1MC�Ǆ����B�a����̦�Pr����gR>���@U����cc{P�N�����B�qA���<�;cexԥ���Æ{�x�J�sV:؟U������1nj��T�<m˲Ww�W{>�HǸ/��y�*�������D4�ȁ�;����E�S�W�PFۘ����D���mH%��p�y��W�f��m��q�򪠗s�06i�@�{��"���Q
oe�n���Jr�7�V 憎�,B"j7����X鐘B�����4�F�DeG_��[�SLb�Qǆ��Rb��ew�N�5�[6S�v!N`) g���f�_��B����	�ڸ������;����y|���i�	�`5!c���r�mH<[5Cn���c�+J �ܻ=�=h���������$#b�0ƹS�4�"�oU���YrAb%�/��W��{*K5q<�q���0m�;A�[Oh��ӹ]k���ކ� �&m<�#s9����;��ٶ�h��-0�mv�"-�}, �����e3Ҥd~P�~^}oo���V�O�p��*d���H?�=׵�,�B��X���S��A"��a@�y�"�� g?���UR;	j��M.P �X� i !Ʀ�4{�e��\�2�<���1���!)Wh���Ls�ָ
�]�i'�H8�M�|J�rI�y�?��߮�py�h�E���]�f���O^��t]}$)�r��郪EdPQ����7��3�1cN_���6�ɧLS� vETq���)�sWq���Ҥ��o�2}+[u���L�?/F��.���n�3�h�TE5��������&#�-{+I�Ӆ:2}��h�	�w}������56?���ۏ)H��]��N��Kr��y�����裇y�볭�>:Pf�b���<�U�3y?�5ȣ�i����p���.��OJl�})���a�3<�8��-�vmv�'/=����SP�^*�&�� �h|�Ь�9CkL���"��ä�°���:֤����L��������d1/��Y_��FYB��0�~ɣ3	�>��s�Ʈ��r������d��'��ys�_�k��^��|@ذ�;'�6��������}ub-
�K!Э�J[h�wE;�u��.��㻷�;�pS��%�I�|�f��فgt+$��k'�9wg��[-������e�3b:����G�cb�b����o���¨1��>"���1��pg�4����J����X"���<�'n�x0�r�����Ť���+�:�[wn)~�Q�r�"����A�U`�G�p��/B��^����������G��ڨ*����#�&��*���(�
�	�p��c;�W(�߆��5�ǫ^�D��@�����Y��O��w��J�Y�n�ÉN1�8�Y=�Y�܀��a�I���S���l�:��Qxk�x���K!�c��2�9f��qJ<��� ��J-Nq`�T�(Fw�#]=ϕ�$J�I��2�Y��f����Eh2�D�YB��܀ځ��ܭ0_��N5�Y[ߤ��,��!?�K�s�#��Zʋ����14ƿn߂���D��d���E�n��и뽲��4���S$H�r�^��j�`+����Z�\�D���l3 �Y���Ƨ���֤*i��'ڗ�>
@Y�A�%J��4�R�%� �6\�bʓ�k&�Z�&�r{���*���b��+*m�s��\o�n����rە�f�����Z�)���kc �N����&j�0O`G������������A5x�z��e|�n؈u/�q%��cz�Ŭ��r �yM��I��j�h�������jO�v ��8�)ز�H5ǤK��z.t�;;�J����m��dK�� �u����d�b��d����H�:��kx�M���8b�Whf��G�I�d�l����o;�e��w���J��Y��0�( S?����l��Gm~����F1������]�y�>H*<Z8�^�$�V��}!m^oW�Y���Y�r7�o�_!m��4yaW�ΰ���Z*P���8�J�xS%��J���Q�[D��p��2�!<�C'���<Ef2�f��d���徝'�Ί�W�a4.��I���Y��v�� "�W~�q[�:O��$;��iA�>i]s����k�D�o<#�=�k��r	�ZoR���[���93i!�aw@;r|�wR������Q�+<ZvE��/�c��O#�i��uϥ��U��f�q
P�m�����d1�-?z1N�^�]�j*r&�z�t�ܩ)D`�y%"��;u��Z>?�����u^wĬ��t
l�ɮ��Nev��}`5$�;е�\��Wl�� ߌ7	������s Ԑ[��q`��3J�R@i�u�Q�����@J�-ʖ9�r	uN|f֙^c�9SC�EY�����%iڥNq��5�Ǘ��2�]�n���nÐ�>y��o0�zǢta����������%�Z�)��UH�Yգt4;#x�|���|���˕Se\�O�����4����m���A)�k/�X����,#E�X�6�-8���Ɠ��㤣�V��4c�J^Ur��0mZ��Hq�ɝ�(w��4x{ϷN�0���q`�n�vgQ���:�C��m�1m� �� L1 �R�ߣ��N�g7ʣ�����rcP��_��~�Q����W�*j�iԨ*����2A�����ye-^������d�׺����|�AE��=����@�<oϛEY��m8�I���\`�����9L�|������8���2����B�Ϟ�mCN_T� �w��g@��n�b��-=�F[y� �����X���X���
��n%I؀���x�����̷��mZ�l1���]�V�]}�غ1���/�7�`���q��������aq�fL�)i��/��?8���j��m�j	�%�_}�F�>��=���/���� %��ٞ���|��z�{�%��,�鑩�М�,1���(\#rz=/A�Ȉ
%g���p�� �����U�i�
o0�.�h\X�8�֋#��qP��5�_�ii[�V���僙���W%�C��m&�+�>'˰�27�5��C�OA��`Q14s����o�n�ŝ1�����"��]��-?H);<�Xz�YkØ�Rׯ��C'�|��������S�`bE�� q�Y�1��e!�{	��ЮåqO���(e��g��������KܬW��9�(������R��>��<-�� ;��Z�� y���^��1[]����{g��xgų)	��Tσ1oZy0�N�n��N��V3\�}	�[����ӓ��|���YT�)��{��Ւ!�t[�d����X��7��u.�V��^��«ZZ8:7.t�Q�
�YnE�ʩQx�t;�%XP;*B�m�эt:	�Ӈ���$�������Ͱr7�p�K*A�v�<D�ÙR�C�4u��**6(��U�W��)������T9�ՠ����EK����$� #�ͅ�����k�*��r���W]�y�0�匙�*�l�1Q�p��
��|�;kA%nC�4Tq�J�kЭ�C�*��7'o��T�s���W�$�#G
y���I:%e8ͽ�8���Pu,/�}���k����$�jm�o�rw��H<��Lb�N�Ac���)�ܑ��ZV5(��t"��ۢ3"6���3z���M_>0#�2E�m�"C>�w���k�"�0NP>��'G.}GR�s��PQ7��K�,��K �b�~�;�B�n�^��T �p<��P����K$�2��	�3Ϲ?�p�%M�l��J���;!�N+���7lGӉ0��ǍD����z�'6jFG�⌲�B�\ؗ(�|�;������:/�b��C�fY����o��$���k�%h�<��q���wQ+���Ю��^z�?_A��tH.'���2\�+9g�p5σ�b�N��sY0�ʦY5h/�ʈ�Ƈ�C��#�;E�����QV�'Z�6�ő�rc�+��4���.� ��~�3��'�I�y���jcRBߒ��Ʊ�e�g{e��g�%#��l���¤^�R��DV�����^��[�P�I�C�xɣ����d#��=������jfd�V��'��^�y�rw�<��
��Ũ���YNI����o`f'���|�y࿌�QX_ǝS+_+1�Yon���Mi�<A�(�c�|��������?55;`	�j)�N1?�0�l�AscO��/�<��H��$���N���/[�Z�a~�ٛ�m���l��
~�����7����[K_2����\�xU�r$�lV�~ec3_�?��mi�2)�QW�vX1}K}藙X���Ń<�٫M;�g����R�)l+���/��������Gn&"a|�B!��8�1
�eNסG��.��	����o�ô���'V��P���L�o=l�H��ڌ�Rc�I������7�#���*&3��;��d��1�3��B���X�7O.<qo�V7s5��^bS������B��gh���8�m͵�^w�&ԭ _���'�B�K��O6�f���(Ǽ�����HE;���<�(��qv+6�u��A�3��D.*�B����Z9_ޢ�:h,��&u���!�7��U7�F����1�a}�� K|i���{���}��U���O$Х(˗�x����a���S����6(�io܈Y�i'�bfG9�� ��f8mI�҆:�T)媌xPΊ��������eQC@_���DL���\u��@޳m�ܿ��&F�5X����?���S�M�4X}Jz�����r傲��_�[<Nǒ�Y���QX�9��v���qG8����+�g	�L =ږf�y�b�^�{�d�4V;��<��W1.Z��^4�#���0�5.ir����ӽ
��[7��u��l��f�ۄ�����}�SA@k�A),�vmE����H0����mj^Yv8IH��G�D9�7n:$��iƆF�JJ�r��t�@KH�A��}�(�TV����v�����7�+���U_�'{���uj!�?�����c{6�=)��z���_���Q�X�� T@��y�Ն�++_	�Ȑ��P������hۂS����xљmf[m��W'�g[����������n�2��D����T��`0f�ҍ�V�\k0�F���0�:>�c��Ԇ]Τ��cU������4��Q��`���I�wȃE�Q�м%A}|���O;�X�i�c��̀� qNkB08��%�:<5�z��1������n+�t��h͐
�23v��KGE섖q�@�wĮ]��M���řN+����.M��������Ο�gc��$?d|�"0�ҥ��_��Ѻ,e�^�=��u�_+:U=%ٶ��?��3��X��C;�����-�CH,n����~�.EC�7?�;GA^�s��Z�ߓ��nԴv�w�I'�A�t�Y8��<ǝ3�H�����)�px���
w�K�.����+76�t�x�u3��8㲚�l�K�dAD����Μ���v�d�YɜD�k��}�e�-�J�j�7����F�BC�ĳ!Y���U��'���=��B3He�"��P�ZY��EE��p$�`G�/���>�p��*�G���%���U�u>��g����j4�6�Ǒ8�wm��./bd��o�u17������QM,t��#�yd|��<��~�i�[�>����h�7\_�*�J����4�7̀�x����N�:����[��\�'���,�j���+�Pf-���*	ޙ��]� ��$�?!)J�n�L�il��3�aM��N�X[~_?�ъ��Ǹ[:H}!��r����e�m扫�{�n��e^Eq.E�Jq�����rњhUG���{#��z�2�7�,����J�xO� /M4ihV2���]��mڷ�Px�H� )��"!���Cj_�ѡa��	�ѮQI>ɡ���#h����"��fV������E5���|�M��, �Al���Ez+˘-y����A2����98a0�.%�Z>�O�y���s�twI������=`U3Ϊ�7�*j ��T�-;�%^G7s诶�,�/}Y���'h��*"�ۙ#YՒ��8���+��U�ځ*с��Z��Fꨆ.�n�{v�w�z��[��C��.Cw��>c-D��@�x�qv�N�=e���D�=451iD?��d�P���n��糩gA��8�>��/�z�����@���$����e!bO�����I���54�@�A���TY� IM�2~�$%�}I�e������~�����g)�I�+[U=�81S	���#�p������j�:�Z���fr������kZ��r#K[`s<����ʕ �Io���� *�ӰjJ1$�^��8������P�u��˭��TI��O�b<��:��L"��8���+�r�,���쿋ԩ��@�{cJ��Nui1S�6��}����Cᴍm���(V��}�s��#I��V���ЛϪ�T
�6�KK�4�[r$���`;�L��N;���ԛ�[�/#K�ix2�j���	m�L��]d��_ �ͽԥ���=�QY`~�)D���Ri�ζ�c�]�Y�L�=!�Q��=��,��&=U�\q�>su��
�M�Tu��E�0��8�^��H��9�U����|):�ET�=y1u
��H�(}
�_�i�a��e?�ϭ�j'!N�+"���w~�A��e^s<Eľ�7���=�0�<��Ŋ�f�O9c�(�FYL?���`������7���_N2�S䏟�i?��Jm9��>d���\<�a�m���pPK�*��9E� A��RZ��ů��G��ó�R�tpKrT`
����If���mY>熥�oc1�k�!�a����#�4@�H�S���*\�q6�U`�<$Y6c�@��"y�D���8�	�@���C�I�#lV���7pjS� 㶵D�Ug��a~�A�,"��I���FXT�Ev4�f�ob	�4���0��zm�ֽ	j6"%}x�������Gn,���8�-�/�� ��_�:�K��.sD�>�O�5ƥ �Ԧ�<ђZG�lk �e{��S����p��4w�4{|�L�c螝�7����tV��߃&�0J(�#膓5Te�q�9g|`b[z�V@a0h�4��s����f)_��I%�� �Q�Zyn�
���62���H◇���y�X�xS:��9vCk���5�e��Gn�v7�!��4s�<��$[��59�f��m���e"ૃ�-���y]#g�����6�O�z�M5t�Ll6�����;�Y�Zu"0��lDa�Ԣ��"���<H]��}*B.����\��<o�ʝ��*�(f
� E�d$3��|nG�e�W&B��m���i.�@&}m�*���%�g��P���"�= 0h@͇�8���b�v��MeM���u�;�?s�yK*�T�,��.u��C����X�M^Nc�!hf����~7��K��b�!�H�Wed[W���o�E}kg���lo ^���q$d���tpE`�'���I-x��+�}���{)	���/��W�>8���<
�~�����s�R �?6��0Q���#��0m�P�@��KZ1�}���o�a���tb���Ud�R�t~�P����CبM̈́���L�]�����؞.ȅ��;W��X�����.6�|�1UZ�z7v�~v��>����+2@{�|�&f�W�^��!���*��1F=%��`P���%w�x#Rm��ҍs�C�X)��z
���or�V2�����)�]I�$ɹB>Z�M�IH�w���DQ�*Q�a�!��#i�[��̀V�B��w�/�2��x05���:����������<�s��ʋ�;ۀ�{�6]�W _�8c{W���"}|H��̫Y�#I��|�>��;l �#d���*��0sV�sC�N�<�+��9�.��n?��&K�����uHɚ"�O���/����*�[ȕI�W���b��7}�K�S��N��\�-,b@­z��RYY������ZZe��M�j����7ⴣf	�4��;K�}��*�|׏�z����C36{�0��/Svre<4��C��T@�N���co달zuD���7���~�it�	GWe�#��Ѫǖ��>�SZN�5��x��5���r��MöK�И�GL���,�y�7㊡N
�dJ�ѓ�Ok"�Y�5�$J{�)�67�"�U�  ̽yj�f<f���B�E�f�th|@���+�n ,�Cupɛ�N�|��ؔN���1�YE2f��k�'o���ר�����C�MӾ��g���/A�~��:�l ��,���2Ҏ���RP�U����V8�q��P�2Ȉ:IaN*���y�o�/���������.���UQ�����5_��B|,�X�<��&�{
y�c)fK���-��t�A�B o�
��k�yH�^���;!��H��ov��|�@*�kݙ,�i�M���R��q���!sP�5Pv��+ՕMjQ�x��`�h��c]DIa�ߏÓ�	��Z�����r����ղ43�屨���z/t�<�=1}�@8���8�����2CH�N�����u蒳�4 �Dc��C��_��1(;����� L�����m�Ĥ׶����D�J(�X=dU�T�v�/����O6A�3e�
�k�f9�/� ^�B�0�x7����=ؤ�-�R���)��������8�پu_ǃ�5�aT�;6	sX�{� m�����XQ�nV������]��P ! ��^��d~a�ܔ)���m��&D��s왟)a��嶺+@�g� �;Pz�K�|�j�L�Rt�Iq�����A��ط20�8
%e��m俅:��-�j�)�&̸��b5aprxi�zI�3�˟��	>��������zh&���k�9�#�ʝ�����tN|�<�*;�-�
�7�Խ�f�:%�4�>w<�lq��x��`���1�r.j�$˖��h��v}�TU���*M��ƪ�����G���,nG�ZO�J��<A��m��p��j�X�sU���t��I�7��7����gۼ"l�$����+(g�h�)�ֱ�f�O�G-���'����MF����R����&m:fV_ݢK��1F̞E�W}P�?T�DN�+(��_*U*r�d.iܝ>�h|U��J��(����*5�K�9$g6��k�4��Ϋ�EΒ�~���O`t[�KkΌ�f9z*{W��IU�΄��|��\!������ܨy2�s&䯂�W�|+Z��]���+��p�@�ۦ��]����mF�_���S��竺�k��E;�����N7c7��z������ n��=s� VA23Y�6@�q13hwQi�/�H�J�9��|�����Q���NP������ޱ������9F��n�fM�,����	���Z�N�S�4'� ����C|b��Im��kc҃����| ��&R�'>#�b���^�Wlh�5�V�xw����L���^Vr������qzkh0
-���
n�,Rw�#ژ핎���u�}]�)bǌ��A�dLV�k/0#~+�P�t��������n���)e�V��qQE�!�	��Z�ߑ�����%i��O���ӡ�T�G����R�^Ϟ�y���~������*��(���]��<$qk���:��*F
��;M����8W�؃�51U<l� D�2ݭ�^�}K�z ɔ�ߊX@.{�9/b�NƬ��Y<�b.��t��t1��6��lA��+�W'�~�ݜ�&
�ȋ���ĜT̼`�x��N��L>������'"�t@�'����T�5b�W����7��^���|Dg��+eŢy���M@��ր7o�Am���*0 j��ѳŴA�,�6�?���Rր={�H�:j4 �`�R��8)��9��(}�v���R���U{����9���b�[f+g(���8ߴW�?��gX�D�0:�?^�/n,�p�������	oD&7qbw@�.���c2T�Yh+���G�Cx�@%^h^��'��y�2g��V;�></�����������V1WZ���t����:�&��4j � �,NK�a�զ�����M���湱�=RP�@���� |���aJU*�����B������_�w�9l�����y|��S5�����
�ǣG
,�?�T�kl<J���ta,t�ڰ��Y,�ޓ[�yg��*��C��w���xo���ej�V�՗���~�������_0?��"��(�f<5�]x�m��˜MED�U�Q��s^J�:�i-E�˫=��f������������/�I-�&�4�i�W㡷Gm�39i~@VF(}�4�yn���6�w�q��)X�GDl���OR��sx[K�\-k%�:.o�,!Ԡ2n\�]!���o��J�r�R�<��H���/HE��`ft�zeK�l���6`��1���Yta�X�~����|�"E�K�ef���'����"�Ҁ���s��<�8P�����Ή��G�Hbd�
��|�6�7�&Bb�d���� }�܆9����{T5�N��Gc^y~f*��v��>��e����>c�N�Z�/��פ�**C�lL拉�'��&��,��DwL��N��^-R{�k�甆��k&4~䆿bvI���*L�J�bi�����!	��e�����A{d[�@_�%9?�)͎	�x�-�vġ�Jk��%�U${C�G`�,�O�4?6�E_4�+�9�����x��o���+Aw�G=+���Z�[�迭tH�1�-s���2z��z�SA���u)Y���U�C��w�p��]����>��zp,2���=�2v|�Q��0��}���"�y���_8�n�^�-7)����}�U2�7��od5�6�+��|���6���c\W��ٵX���B�*����]���Rt��۩B�Gޟ�����6�}�5{��gե���^������)�*9�h�
��O��g_j��Cv����!�Sjk����f��N��l��;�pI*ʙ+���{��|��K�[�b��p<JE�Ժ�p���=�lQ�)�(��|L4�N\%d.$@�8R�%����~��N�yJ��]c�J��1��,�F�q��|\戸�_�*��o'�L�܀�3��l���F�ǣ�D��9���d{�c���u�e�l������ؘ/�F���A��SA��	�Z��q$uF;2�<�/��q�hJ��J/�J�+�5�#�R~�Qf�L���0y���O�SG���E`� !����]�u�����7߈��B.�B�,�zǟ�����&������|� �Yv]R��O�g��^��ٜ�O �e��TU#�lq��7�D�"�����=��#�&W�q2���:��4�a݃$/q�kFVs�#7������7��b�H�Ep���LU�:��G���[�G���n�4h��3�+�����1d��6�� ���/ANv6p��G��@�^#/j���2�z�+����	��\|�k=o�h~�݌���þ��1(t�>�%�s�RXB��`5��<�*N\������m1�=u��k�r,���a�mc(r��Q5Mx`N��ߖ&>l����el�_|_�X�y��H����~�6�
��A���� �3T�lw@-��1V��Իv���k�S��NLA��p�����c���+f��3\;Ha�E#���|g��y2+5l!
Pc��(#�*iX�ɨ�w+����l��/�H�A�����;�"��0��S�7(����(�E�%�T(��$Y�c$�_)@�������bu#�x�@���S�!n㫥�L^n[���x�Y��kf��L��l�;��C��bmP4c��gYy�o�@d�4(�Zr�W�RJ�E������8Ξ;�G|fG���t�qRB��K���L�Fm)��s��j�y;Lb&�в᛺DfGqHs-*r|<�P�����G<��2R
�3y�D\B�J�?�����dE'�B��)a�m�\�����$k�Q�5�(N�d��80���;M�w�UT=�29���<��Bq���6fl�_wԹ�*�b����k�J>��kkב�b��n��#A�z��dl�S�v��XWjNpvך��b=\#f��������$����|�Gr��蚊+�����X�l�ˠ>mY��������_8I/� ]u�e��,���q��-��0�D���9�zŷ��S���*�9�C�'|�t��em����m) ��iB̨=�
�'.v�=	i(9�(�5�ƾ��Vz�K���y%�����tq��#�6���%�&�E�ZuڭNńz��(gw��l��1��`��
�m�u��J���Z&������εu��K�5+�4��$N��^�Y�L�"���_��9��b�s�;�Z��pr,l��@����.�����ä�3DM�dfG=��ؔ�$K78�䥗�H��dB��V�'���W|���}���'h�w>̳�urS՞\w��Ww��np�צ���)K�c�BLDܹT�SO�^����