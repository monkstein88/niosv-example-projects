��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2i�>�|���B��,<��\ ��W�~��O�?��K��<$џ_�!�ʙ�E��7<�}V���O�~��f.n��vջ��u�ֽ�9Q�>Gg�|�إ�ښ�9�>���r���_?�byw�4����Jn��ŧkg��F�<u�U.SX��t�K�h$��I�
!�{��<�� ���$�n�_� ,�v�9��ft��̴�*&%�s����x-���](g�3�ύ��S.Bjػ%��r�l�,"�a&[�����mװ����6rP\��|K������9h�?p>H�1u$��฼#��@����� ��f3tՆ[4h�ͨh�������a��kT�x� ��	���#���@��7t�d�/�S
���9�I% �!���{8'D3X�2��J��/���ϋV	�lYZz��JS�� ���w�m�\&`��0Ak��H@��7y��o���V�V[0>�����(a�pxn˂\E0Ԁ�p1?t�7�K�h���f���Bn�KC+[�;��]9@�Ee�^�t����Y��`�Ni��/o���ױU�FU��E���o�%T��9��7�rz��wK�Ь�=��N�A�:�R�r���Q��z�i{����>Vn7�U��V-��R%�Q�R��e��}�����z|ʛD���b�v��d�#)��ţ@���sE[¿�D��䂓5���>\����;&[��Q�/`�.5P��4�OM]�<3�@���u�ל���D� ;JU-�F����\�}�6�w�� �<W<�kN�C��Ƅ/�Z5��^,����x�Cw���O������7��h�mB�I_7�M�v����bQ{,�C륳����ي!IfB�i0�*��r�,�AD@���[2o�����7-zߜ2��PjxfT�Y�w3�s�Z	��C<YW��]�!p�I�����^3c1����֐Ιz{��J.s��U �yEfqN��(qG�	���gz>���ѕfv���ڎu�7���L.����zH������ɐ���-޼Q4 ��Q���
��cV���!Q.��~���s����%��k/T�!���ŞB]��)<'��#�>�ѱ|�\Q�R����zb vѝ��V���,���u��Qp)���*���\�	�@�휪�49Lbe���R��]O�P���K������@�X)u��]�a����+mt���� ��aі��
 '�[�	vH�h�f(�U	U�L e������a����(�<�a��%)��M�H6`Y/#���2pPa9�A��������Td�*�ڤ��3��n�-a��®`�\[3I8�3by�`���������Qh�ҕ��fY �7�de�s38���E���:�k��	�x}	�'�`��� ]ܥU�
L|A�2����.��Z�z�Z�n��p��7̏Bw �'.��`����gU�S�G��6N�m�N{��+M�?��	�InL� "kH9���~�m���2�����f�,Q;4;��6E'�1�R?�W(O�r#�<7A�t@č�Ѷ�mQ�]���y��S�("i%������eY�{ep9<G�y�s��������^e�aaN��7MJ�U���ӯ�_���y��䑄�Z�5ί� J &�w����wm==���Tx%�B�Cln�pc�Z<�(�'E�	B���?��� ;.R��vS�Q]t�cD�=a8�s?�J�m����Q*Q���&�Z[.&�v�)��ʚ1Mȣ)n{����O�IK_�/��B�@��Y��UQ���#��2�PvQ-���倫I%��l�����g�����,�m�/Z�_��x�ӂ�;ޑZ�6��g��ѡ��0���l�$�։=[�m��&g)�R�Nw>�oZEVݒn�e�e�*Rx�<�1��짱��|7��k!���6��
2RMpF��Ēw��W��]1�"�l��V>�x��h��`#��3�ƪ����%?��"���+���YJ��G�-�8�Ƒ�W�
�XE�r�Of���u��g`��R��Y+��r֟4Ȯ��,�<<�G���*���ʕqX6�j{��ۋ��Pw�˴�|d� krˁ�� �� ���(a�	��`o#�G,!�o-fi'���$'��$��5Jr��O}'����m�J�+' ?D� $c�_l��/�"FF���=k@�(r˗?�u�s�۵@Ʒ�	bx-6IN���I6�\���s����nxM��	�D�p>�A\R�� ��ɿ�T����߆��*������������n���#������m��A~��?X�B��Άj�Z���8#�Sc-�y<��Y��O�gyJI�wx��7�VN�	�wDY�5q��nffmk�uW��wI�{�M�?�ݴ�����t�|�Aw����s���"��,��6���2�E6h �ғ�p{��!x��;�EV-*�AL��G��r���`k����Fc��g����?�i�U��!���y��~��sq���B�V���Y���CA���&Zf��9�ʉt-?�m��~7��L�K��Ԧ%�mN�y�Nw��!�I����F;">�M k�t�6�%�~����VF"���
��xk+	`�D���KY�c@�v����Xi����3����U԰J�>�p��KʹU ����B��B�í^������G!�M�I����m����`m�>.B��P��7[�ߚ��	Ge������H���F��N�IP������mG$9�f�����S���
�2��_�Y	*�R�W�)kIC���Qn�����Kߜh��)��G��V��h.�T�:߫�����%���`L"\�y�t4�TC;��7��BR�w:�yV�BB���@){*�>w�
at|Nmg�C����d�"1�j��[�~��; {�����x�Y�5xᐈ �o��5s۳�`�E�i�= �]�.=�B�ûӅ��i�N�J��)b���$��!%K�̛ �O��e�6�-��Z��������؆;�T�Y�s�1 !("d�C�lG;~3�nO���~r$~�9RC<�-�&w~���6��˚l���E�'y���S�:�ƾ��N�Ϣ�kQ����c�0�����&p%��h��C���)�����e��il:o�;[�e�X�H�=b-ϩ�\/��&8Q򋿒�4��n�or��OWC�4N���Jߛ�2X�������J2��)����:���~bT.^���`�h��y�6��m��➩��v�QMȓdH]J(�LX�z2��Ϯ ���bP�L��X�]�Ș�+p�C(���q1dD����=M��*�aη?f w���9�"�wԛj'�{��L5�H6��(����	@�����p7`�����t��k��>��)�	9V��j�fz�1Ҽ�u���U`�@P�yT׽p���~���G�Ç���`��V+8�7wy;zn�sW��|�I��,���ĊW߫�� �|ay;,��*���?N��}����S�t��G���W�a��(�ȇ��F82�\Y��c�K6����n��.L���kQZz��:_�״�1���J-gj�_��k����yd��\���9�?����%"[j��Z��~��v�R&K���E��q@�F�`>�v
�j\�Rg�,7�E(k�mk�R1f�P�
���^�<	xO�VwƂH��$:�PbA*��:ݺ�E:�5&��\eq�`���X��r���j��%K�"�d�rs�g}E��ۿ��:���}��ጆ�{�g��4F�������^z@���0똅,f{�B�ܝC�4��"�m���HJ	U6'�UF���ψ�i�"�uY�?a�_S0X�R=m���Od)���(Z,�w$r�c���f�κ��b�V���S�<:0<��$�_�p�Y[S�"�nj�>\H�]����?ü��h0^�~ݜ���9��&��T�;xpy;*�x��Gʮ9��)/-��N��e��^i�v��;$�N��Ie��p�� t��O��>n��[���b���#��X��E��1"���#�A�ʳ���E-?{���~��d�tҸB�8�����;�K��pM��4_�6������MYQl*p�B�+����]!$S��C�S�� ��=I�6|ӟ�y�i��jh��n�-;�NU��<nC�5�<H�ՋM�z��g����9���K\�����3���5;<2A:���e-�@�z@hQy:j�Z��J*�� %¬�b"\
�7�Ԫ
���;�!�_�z|�y���"	�@}�բf/!Н�i�Җ�ϕO��C$�Wj(���+�A��a��e�ze��<�5��A�*�=c���6GL�=�&��
�	(
��B�\4ȣ��w�	��K���b]��b_H>P�*���9��O���l�v��4��R6!�"=�3[H�:U�A�c���6[Ԕ=���UI�u�e�(��j���jG�L�9��L_��߂��C��F �HR$��l�#W�i�b��5����ϓE���!Lv"�;�H�f��u�s�"}3�1�(p�So���?A�[����SQ��3_�|B���F�H��xs6�T�q�
C_�\s�fuV�TQ�_��I���%��k�����߮�v;1{��hcc9���+��o;:�윇A!�4	��cZ��dI��͋�nuXCGYz$X$&������qz+�j�r/b3�a�͜��}e�|�2��&�2a�b����2��k�w L��	�a���
��7۝^�Fo�]Ԃ�m�JQWXz��]ixqM��g*�`��V�D&*�2{�]�H�@�:�R�@Ng���S�z���D�iA�>��u:�4��cn��)01W%����oW�;D\�(�IYR�ؒc���G����qXrd5f)-H�����~eyJ��K���8�/{�{g��KY�-�ܐ:����7O������Wm|��u����a2h[b���z�0T���2�ӥG�G	���՟�8��i}E^hh�3o-r�S򿮀��1�ڭxnd6�s��P^\c�CFg�������1��,�)�& >-��5��(����	��/h셾�p��L��9ށ��h��1�ZZ�6)$O����$��+s�lb�C@}�%��I�.Ub�05��@Ѐr ���<v{��Z�풖s��?<��N�|�s�e��^��]�3��>1��������|ԜGZe� ˛v�R�>�K�"��� %�D�����u�@�r�m�ȟ0�; �{��3�J8"��sS0��}�_�Sʽl��+���S"HNɼ�
ǅ�#h)��q�*�%/����9�L/3��`K�Ϛ�H�Lr���X�W<�1	�jܯ r�`�C0o4HX�}�4��M��t\�����VL3��ƙ�|⊞eُ<t��5�ޫ�l�X0ce����Fz�<�����ڳ3��ս'O���0��"�[,���r�/Q�@_EaR`S�ٯ�h���zYͦ"V�<Ȁ�]���E��Ӂ�XoQ�� Q�<W #��ً��H���|�7~��;-�\�B�-=�� �