��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��0Ǟ���:�i�2����F��Cp�٧�%�VU��^�}���wWN#�|h2+2D7�ҸQ!��,��Y���h3Ã��]�
#�۽}�0��TUTE���x0#m�k%4CxK���Z��p �k>��s�G V�JuNGP'E1�f��urW�;�s>Q���ER˨�h��%GNr+����5�N�ԛO�3�W��N�'�e�.~�a���ݟjr5��T�}���s62~|__�>U(�_����S�?�_�q>�]��(0-{S�Y�s�6Tp��mR�C�L.�T�b�|���[��2�3��L���j�U�⣃^� 7I8��)��;eSpR���G�NOA�sD[
%��<\A����Ya-;�]`���	M.S9kʾg�⮀�9P���g��EQeϹe���%��2	/�lˤ`ss �ED�ǖyk��C�lҞ\7:�p���h����2αc�6�1�Pȏ&U����U����S�q������ ��	avO��ʈ
��k���Z7])Cv+����3,=����3�`��Q(n:8CG�p�Z�V`C�kw��[5�R�6o.�Y����a~딃S��c@��(�v��f74���������y;�Ə�"]�q5s��a�zί�'\����ڜ��NΈ��B�g26�3Ԡv���T�}��q�f��h�QAO�>���b#����xi��]���Sh"Os��:�g����@!�6�=�!���w�����De��]R�/�G�Nu�˅��i5���Nt��Ǔ�65?s�|э��%Ν^(:�εp�O=���*�E5J��3�@w>m_�W��QB�j�7۷�睫��F9�ڨZAK���=<�����Lb����I[���4��	=��7���ߥ�܂�j&��
-F��U|)�����T�r��U���%���z_��sAF�a��P���dR;2����RqJ�XJ�^X�������j񳱐������I��u��Tu�y9�oܣ�f]2�S(����.3à�܎�������ވ���QL��?��}@�ohv�i�
�N9g���*ϴ��
������|�7҅�Pv8{V��L��X���K��I��kG�r�G.�zU�����Q~�5�FT��u�u��v�:���f4�o��
d+�-h���� P�k>�����7�l�����p�CU��a�mX/H��s<Y��\�t
Ne�F('O�U|��ע{� �����n�oI�l�f�8#-�a���
�9���ĲDv�P����]^�%�MrJu�MA���7pdx-���]��Jp��}X�����u
^���tЕf�Q���Xb�\gW�x���ԁ�Ǚ(xQeK)��>e[3��Z���T�=����"䄄�u�8
������~Gwb��?j�ļ���$PR��t.��Rݩ�B��y�rg/c�:k�V� �8��ko:�	��w���N�.�q��f�P:	bHCb�в�6� ��w������������P����Î�~���)�բ�.h������:]��*���ɽh��S��&����"�"�&�t��d�k5#����w���24@(S�S�'����
�.�]�,����dđ��n�ұב�4�Z%șBx;���JO,qb�� |�ǺĮ��W%�Px��s�(φ�#�ݱ�O��B.�vz(�5Рg����±���D��Z)�zt�吒���Z���N��Ǧ6�D�X?Oy�d.	3�kJE�C����5��ѳ͕���h��H�Y]%�	���J%�S��q�x����APl��E�R�(Ǎ�����Y�h���R��5������iWW>��7�E`�u���٢ɴKv�po�ӅD:d�)�Zk)ѐ�bEK��)''��z�S?�����C�iX2�}H����/�Z�zU��ICq8�D�!,����WD��HW+ ��.����.Ũ�C�l���<[9��V����	�#���X�M���Rm��6�^�,�3`d@
[a�oIW�Δz(��CK9~4�N�]U��Q�"�GY�ܬ} q��#��0.�m�E�ݦyv?OdzS�=��jz� �I[����x�)�|��|7<�~&�R<D7��G/r&�����mt'�܌o�,�9�~W͚���l��,e����{;��VbQ�ՖŨ�fDd׹��Q����'d�� ��we��h�0Wz�]K5�SE��:1�V��{n+���_�CϬO�aL�Ra=�zP>���������~p��t��I�F��j-���B��0�q�Bz�����H�JM6zoj��uuQV�"�79]؝�b�#d����rI�5�iܮ�~���gi�@|=|A@������G��yA"�b����q�M8��Ą�}���l��1�˸���B�� N���<����6�p����r���>�+t�C;G�6���r���V-t��T<�l+W��Ak��a�^�΄��C2x����TK]��9[�F�_%�A�F?�P��ȁ,0�U���K� �w0���������{�t⇨��l��֒6���J��W�*_�d�l�O=�Ȯ��/^F�qC4�Nk+}.�2�
n��(?�Q��X������t\K�J?��%䎈!�&LӼ,�뤙#�H��g��g�e���s0��z��^���d�Zl��Ź�Jx��(�i��5�	9���P%���<M�+���o��H�R �j�O$����l����rI �'����Ż�]<��z~�zZW+�+�`W����.����TRi����%LH�	t��Li~L3V�e�U�J&�DUJ���~��դ�������a��=��aĤwnF���a
�ɰī�(�7v���.�|߷�����)>���i�v�ڐ|^��*��)�>9@&���"��JB�W�<;>�������l�����e�*�#�S��lc�<��R֩)�=uM[n���xԂ�h���V����a$R�<�U���t*~��8F�`8�,�'�㑗������q	"�?`������xy�U�mm�Df��.�hXz(���z�hu�)��K��.��1����wA������缴�<B���
��h|��_�2o�H���l��gG��=yYU?3<�Ԗ-XD�-��C��{���ê�
�3at]����YR(��\R!��Z|ǁ(��<K�*�m¾�w��r��FgьEW��F�e����Ȩ=�T���ɵ�'[&<�_��Y5��W�%�m�q�U�|��mIO���ٕ�̈B�1��6�
t�g�4�;c��.	E���J�KJm�|J,��.Mmy��W�V�wyO���T����縃�8��}{3�]
�դ����M� ����`[��%�XX1τ��<��|�o��M�"��)s��A���(xGo��@QS7��'d�g_�q��3����<����It�v�ǁK����x&ː}�"j�leF{9�y<$�<�Բ:Tt� D�ŋom���#�R��2�d��֯Zt��'U7����-0��L@U��74x���DJ��m�����*�� �<z̵N��|�X�G�EsT�O\�>RQ�s��ػ�>�c�_�\��D �z��Z��%���KN��pwު���I�LyE��BG.=,v@"��WQҏr5=1�l�d��,�Vv����HtOi\��t�Y�֫��߫.��1�63����A�}��C9��I���屮o��*�_�ԓC��s6�bE��"�g�:*�~�!��	�����k��`W��1��㕄�&�9Ti+_Ռsc���4�H����V
L$'d{�zѨ���W<�����#�T�qY�=F�\��U�wc͠���/�����_���`�/Y=�!�^��y�l�yd_9�����&���v]I��A�cűgĂ���U���Y�G�Q{���M�>�}ү�x�� ����5��N� ���N�N���Oj,��1	�;��-4�#E� ����}��������d�M�#
�_���{i\�U��?��L2>;|��ᬢĀa�a��r�-p�T���j&z�vvЧ�w�d�ԥ�3�]ϴ����8��Ng}5�d��ǯCإ�����uCQu#�v�jմA모�h��Uw?�G����W^U���� it�Q�GI�C�ia:n�Oz=!�8ch�ߑY��5ܷɌc��y$���Kd��!�Q���G�,�л���N^ό�z��i=/¡��g�%EڀiVkc��%�^P���'ܤ;v78X�̶�sƔ�7�ϋ{7K���+�Ţ<%#��<7������n�}�Я(re���@bZ�����i^M.�3��h��>3�C#���K�����WŻ��ʛ��o�}B�_�w�o��	�;GaD1��#�I�����<�����C���V����?d'�}�)�9>F�>�F �9�����_����X��<�4��b�� �^�1��4+������'9\��*�Z���$)x��g��xWo��i���A%6��	E��#��L�SQ!Qu>��m��۴V�9��ՙ	�:#��@^�tͣ~���X�xo����v�'�s����w�;��y�:���ј-5�<���e+���c|6�0�_7�ݑU���b+��#�3X4�)8w=�%�ጐ�
Vҽ3kt7-,I��ԔmDA��I�`~^6��֗>�A恒��Ra'���>ږ4�>+��o���A�	�����'_����h�]�׽؜Q������L��&`���]�E�va?�)関���R�������n����0��^_z�ռh��g��#�����)�f�.oDEw���C���h��@�r��:ܸ�2��
@���^]���Ru]�%5��np��eatX/��ܫ�l&�-*����C���ei��Q��Y�ů2]zF�psF|'�������ζ��[3s��Z��4�ę��GS}�8������8k�)&�.�Je8S��:L���".�0��a���6a_���l��P;/8�mxFs�Z���8��<��9���gd;])˲l����'>�VUt"�=׍fZ4�&$|/��0���>��"��ƶ�t���5䬶�Գ���O��=ܼh"��й�[��YY
�=�%�/��7܎�5�ѝ�#Y7�B����� �O�"�w�
[����V��Q�Ӂ�.�愶Y}[�N0�G3Yq+tL�dz�o�
'�Y�:�Z%E����A��(l'xowMV�?_H~�W��D�`�5�nn	�[�����6"�A�銹OZ���r��	a]<R�O!?Y.P~���lf����"3���>��|�l۪��[V�oo��d��1���
'�	���I��W���ŷ,������Yb�^�v�:�L���g�H����0��7������T, (��\�u|q�[��Ф����<.I:>F���.���2���I�n�!k�����^�ť?��^X� ��oJ���J���$���R��O+[Ƶ�k���=�0Hl�׫�FD���L��:vf ��6�w�Y_�2p�q��Y��r�Q	��;Dh��gȖ��'nP&�`�z�E�C��Es��0+�������kg�2���>�{�w���J})�-�cb����̀�	{d�ͻ���J�nV������L0��(.�
C�|3�rD~=S-ւ�R��0��x� ty����p��L~)���2((�����{����@�/gMQ���@	d�6�+�SX�ܨ.K�t�`���oF\7Y��'�2Ŷ1ȃ�������*�}�8����� �a�����IZ#a>Y=�����3���q��v��R�7Ә	o�z!����~��@����s
tj�!�R����{ax���/��_{�����$�����<�z�h�	�7����TF��Q'�In��;8�6��]�7SyInB��
�����[�HO�|ECֆ(F�O2 Z*� m.8�I\�G)��	��	����W���d*�S@[_���TV��T�|�k�$�{�P�-- �k"�9⾼����L��JV{�1��K��ݵ�_ƀD�X JF�w��錑u�<yJ"�u��ɖN*��G���L�J���r�)�;���\��3����o}��zc0��+*�z��Ւ�)�������`�r�䛜.��e+I��������K�r��J/���N�d��TKRu�2�d��c.3�h�4�`��G �G �����W�c�L`saEMv��-�tZ -y���T���R�t�h� v�cý��������S�v!?��p
X�Ы~���c:h8;�	��V2	�.����tf�f���BQP��}��y����Ʊ��T"-�{��Q-�b �k�h�����6(���4
*2��E3���F-��\ud��4֏�1F�0�� ����Rx��%�?y�f�����alJ�;S���3_�q9�]��G1Z@"Ң�nq���sꨔX��,X�<�1O� ��r�/�ru���ڙ"Бz/z[��(�z�&��"e�^gˑgOYĎ�{^���i ^Tk�~E8P�-´p���:���t�*�7��A��Fܞ��ɷ����� ��J��OX��~��X�m��û�8�񏹢������#O&�aoɯ v�gkKI/L�*�Dy��,P`��5������� I��O)l��ɥ!����������"-{aUj�s[T�<2�z����Q���p�Z/I(��X�z��&R�K�w�����sЫn�R�� �LJ���V�ԲvB�>��ނS>�K�)��� U�D_q�ƃ(�6�q83����P	�����������i�aU���ƪ�+�ƫߑq*��@���M��P�l;S��=b�B�h�T�&����s~�p���p�O��<ͱ���Fm���c�շ�J�K���J嫙)d�Jy��(-��s�h?�5n֞�6���P΋_�O��x�O�C^P��Ot��*��A8N84�`�Z�^�۽��ǃ�+f,Q>ם��Qx�
x��	
�8��^�[�wİ�Rŉw���� ��ϳ�S�!LQe(��m�
�1��f9�%Bs���F��(M�j��_�z9=m^�G���E@�ۑ&i*A���`�`�:��<�U<6DE�S��?kB��/���B����,?����7�J�[G���B<�@���ڬz�^+	�[s"L,�>�8~̑�i�O{� ?:S�y�T���@���Q��$9P>�$r��5�:n3#1%ƭ��J�)O� ��2�������Qr�2}P;k�� %�G�S`�=/~����x�j��yq�\,��cԥ�_K���t�@�´Η��\�����{��q��E'�Yg���'9�#�J�+T?RX4<t��:��A����
F�J"�_WS�	�6Ջ;��㩅�e/�gQ�����38�ayS����p�����f����/I>6��WΡp�w5Z_Jb�RE�� �<Dx�A�ĥPb0���U{�;��{�����-U)�)H�qE�P+���Y�K׺pܹg�W���ݑwV����=��3=����؝����.��k��:Tvj��V3LAI�o�H�]4�Pq��?��8<��tz�8�3���l'�ܦNؚ�E�>E����4'Ѧ��^���\�W�K����S��p7�4+�d�U��098j��X�i�|��lآ	�񾫊C���O]���8��;r
�q�3ө*��-�JlGY��x�Zq�'�l��o�6�J�g*T$�׎8QB�x[��.�3�	WX��z�q���$�+f�\υI�R�_�OtnBA����7&��,3��z��uM�zh)�f�ҼZ۞����<��+˿�cJ�th�ff�|-7�_�fո[��_M���y�2�w:���أ���i�:,̹���ktw�k�mM��Qs%�^�
�(��WV��L\����K��qR��t����5~	}gV$H��Q&vQc�J���(��[�F�LO�'-1O�K����ߕ/Be5N���`#Q��=�j��XܲK�n��8�	᭗����!��T,U�' �Y�di�R����� Bk��}�s���^l�v��#`a�ͩΔ��9N����y͢3��*`����y�dP���T���/Y$��C�lb��XV'�-2yu���� �0/j��-E�����2N#û�k��վ7�|��C��p���H���t��ǭ��q���n�u����SRI��Nr͏Ŕ`�+�㰋��K:�1��*&�
}�c�UKO����Fv��������t�u���qEFj�XNF�g��:�4M���4�m	�}����Q��%k��[ߒ�[}��x�׳�ds����PV%5dG�L�Aj�f�N`H%�O Q��z����?c�<|��EV:�p�� �}���R�.�<B��HEt��7�Ax1�A����L����y!���d �*���(�[?1�]0n��k�]dPm�(s-m��!��J٢&ʁ�<��{G�������0��e�و�B�x��R��=����c����%��XD�F� k�6�� �<� 'R���,����e�aB1.!��4x�=٣���b>��*zךg�W�>=��Bu�m�I��}�\d:Z�"����C�0df��D.Ϊ��&9C^�(|�����ʗ�P����pFi&u���@�=�c��կ}�o����:��]�m)Q�M�@��
��f�)��F��H4U|e��ş��̓.qab箾��Ey�\�Jv�ڡ�+�Y��E�T|���P����`IF�PxӺ�Ra�qZ�эV�W��b���Pʴ�W-]����ؼjQ��5WF��AWNǯm��ZJ.9tRI�+5n���s��_����`�=�|�I>d-UIF��4W�=�7�5e��,���'�\�Xi���N.������� �6���7
j��Q�
﬑�i�A*+e��@��IP7*]�#c�)�y�N��g�$k=�+ֺ�1fDV�����i'����n�(!U�	��E2K��7��	>�%���󙛚�x��5֛;��:�mm�S�3�bKR�;V5 4%�ȓ�)�E����J�IҞ�ixv)�%�������\!;HH>(j�f��C��nk�v�L�P��vɗ)�ۨg(��
J;#`Ě/�N�C]���fr�Z��������AvK}K4j�i���8Xh8�7�a"���E����ִ	����3�/�ȗ� bA1�E%dbVz�p̯�g���,bBS,{v)s6o��U���6���8���/IU��t���)i�W]X���8 ��"nu�de�t%�f��tNT�(m.I�ݯA6|N``���Hޙ-�Nq��n��87��y%�d�],�<��\�'a��L�])�-��{Lv�sS�B�L:H7]���vSa����0�����QU��]��]�*m� >�	�>+�8�1��4�n \J9�W�S9H�x��B���@�� ~LN���k�"*X�mx\NX)�V��B�e%��D%�9WL)jC��$�	=L7fq��Ȩϻ��(�l��]�?ɯ"ڹ�&B����'/���g��B�R��{�d�~���]�	V6F����;�Ũ�	] s>gNZ;��"5��Y��udd��bK�&�R����%�?���|�`hYc9�%I���:2�Xk�n!"?�'L��#*^Uy�dW�l�
L��'���(�{js�[��Bx_	�����t=A;2������ĥF��ƕ��4"�GM��W!e�՞Q�Y!cq��%��)2ÿ��P��č�&�m�+�����d��qD�B��q��){\�c$�����8�k]�����l��P-��ǌ8�8a�Vo��<��� u��F�"�D��� uj���w�9�a��e\�]���=���?`k�)��T^�6\+�5��T�B��K�u��6,�^3���ć�.�5�o���Cfg2���U'	P�q�>��mm�e7�D;�	ZT�������臯P�a��7�%���ш�EݟE�x���c�T��_�x`:�{n:�63"�q"���_��TBߎ�ySLl"-�]�\^Kl�>^�� J��� �
kff$ V�P�	��Ǐ��r�`p�oY	*���u~([���ި�[T����h,j�&��qF+�+Qn61��IUSuv���C���2�|gv����W'�(Xf������ݟ��h�����O���j�\Lu�|�xa�9�,V(�,u��ȱ���{���7=6��x'�+�����A�O��d�M�jzv�O�×��~Pe�9���%�+��MoMߤ)��D}��$-�O�Mm̅����O�M��Q�W����R��S�P�:)��k�{:���Wf��9
<?E�+���������e2��%�5��G�v�J�&/q_��~=��H^����j�OTĳ)$\kr��^�/\CȪ%lNVl���:�������5�-Pb�V	2$Kz��7y;���f�g�J�E�C�^�⶜����M��zj��9L�>U����4Y
p��9���b�nh���\�'C�؊���7P�.Piz�v^�c�lF�2�1���=5�%7�i�EF)����=�]~����4���hP�sū�%��TrV�Of�����U�3Rxg24mngQw����Rt_�Q�C[�%פ�}�5`8���A�G�mh��:�õ=6#S[�1$�J��˭���l�T���\��	�W���u�(OF�Nn=c;���&����,���
��1�&�_� 3` G��:A�_c7�U*'���y�b
�R2��P�6���w��9$�1����-ǈ����³+���g�5�{ԕ�d�xj�j;�L:�j~}��`n
�J;gѐ�Ă-�:m{+�k=wy��}��	�>^�dh;�@G�5C~��poqRE�23�6��s����_4	�E�8&8<���ڻ�P�V%�@^cL'��6��x���?)ˈ�rS_
��?�r@��P�.�+�����7]	�Z������.,xI�!�I5��� �=1��H�[�I�-�q�`@s��.�7�a0|�����C�ً����<S�88n�╂;�<�aR�@wI.��sh�&61Ŀiΰۗ5<O��-��W�r���3�*��ڝ! JK�>��ʏ]`a�c����׶�{�_��L�Kf�s�������̻dg���S�I�@��B���Y�a:lNa2�π�B�	)�T��J���ws�#X��G�ͩ;L꟠�,j`�Y��sd�$@8EǶ���@nx�]�j箱�c��)������64fwbaԈu"@�D�kr=W���?����\a��D�����x�@�/@�c8�V'�;�r�3Ny��𐟶tn������|��9d��)D�k+��:�ٚ��RS�`��P��`�_����Wb�P&P