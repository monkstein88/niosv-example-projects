��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��0Ǟ���:�i�2����F��Cp�٧�%�VU��^�}���wWN#�|h2+2D7�ҸQ!��,%��.8�R'm��lM���(�ų�1OV�k��u����岬4��O��ꮨ��+!uٜ�l���)"������L�r1�z¯f�%m�e�i��qȌɅ_��`G�;?�*�m�?&S)���#�;̆A���4I�KQ%���u�ԙC��v-9�1WY���Z%����Õ��t4M�����~Q)GKdz��q�S�7dt�]mݝ[g8��j�u��`	u�VE� ����&2��M2����	�}}�^��H<5<�h@2��ZUH9�Ǘ�F��.����v*]X�
#% ���K=cN��H����&A2�)��X>:Y'������ĩ��w�W*�S�3�U��:���TECz
��f�>;�ȼ;C�]�Il?CT��J�E�**�@��k�ƒ�"�u�����W\���6��D~��wN��&�\�j��>ϞØ�!��?�D����bٕ'A,}�$N�y��]�e�Q��V��$/&3zw��,3K�<��?�C�gVM6��n��S��Ju�w�����V*��F ���^�Y��H��X���Cʡ@�Ǳ���1��5�ο�EX��E���Q�%�ͥ�b� T�0��^�;+�Ͻ?r���/�U��ɰ�A>���U�1P�;�ok��A��@��TM��U{������-��I���MyQ���|<N y��aH�m�v��r�Q ���a0��`�X�K����j{}t������}&hu
e���pw���j��Ye�� �{��%@��8
�m]T(�1��n������Kisg7%�I�!� a�3�\@�_�B$٢�oY��L�>
P�_k'��-�����C+i��e�!��,�a�}��i`�S��.p�Ef������C��L:CG��>0���K�}Ycq7���3?p�t|��R 6)�+rVi�u�rl$�⼕�O�ĒάB�.�:݆�� ��O�ƅ�M�6�Q����,�X��5�R;��2dH�gVg�*����@��|oʋ۞4��N'��,��wQsr�am�V[����-�����)��u�+�7$���-��( w¥b�_V�����}�GLy6N�Q�zz{�-AR�=������/I��c�2qZT��<��9�,�g�uS1?
9� �;u�ޟ���:v�˘�;#��E�����h��Ag���$g��.���xٸu��sXŕp�{�(�i]$ ���[|R2�Hl�������.�i����"�MG}�u�o�i����}_I5��h3͗�"�u�5 �Q�޽��L��λl1K�%ت��4�1��<��t�E��q�e���&l�S��EvWۧ���l�7����L�������g���XIJ}�/�M6���%�@�b%
8�Q�����:veځ���hrQ��NRv Kh,���ү���MՒ0��T��?�MP�T7�T�j�)�k�Q�T�%�nSW�`��k�C�o ]k�(3T\�W卪+��k�f�[@�P����F�(V];�ZF�ڂ���(�L${��"�X��Q���:���VW��"������Bj�#le�iA�C2�2��Gt�㤬�~���EV��$ĴB+^�g"����ǩ[�vFR��-N��,��A�H���g$��N��v3�m�����u����E��9��]�b���q�k�4���A|u2Bs�$��ܕ�-y�PmDkjϭc&�� �pvo?2��jMYF��hߟ^(���N�g�+��1/L�����9ȟ�:��
�6^�����ts!v��*%d�:�2�$_��>.}�,�q�%��)Zfcͣy�fM>�~'?�]ɜS*�F��7��Q,�C���xh�� ��ÿl����yI����wOx��G�ݵ]�кM�"�͋a^�u�� �Б3��,��:&k�Ժ$3}�n�_֓8*(��T���c	,�	�ny���}�6f$��	�y��� �Ϗ�fĜ:�5�"L�06�I�c����*��R�uȶR��$������w#Ɉ <�D��/'<ޠ��z4fS��3b��P����G�W�j=��X�@
N��<q��>���0��U{?lR7C��Ȣ4�w��5:p���׎+��
�5�:fP����`��RR5zc	#Z�3o
�P� �"��r�B_M9� ��)�+a�O[���8�\k��W����DL������|a�#�w��c�zd���EO���1�V�{�	�i�u�zyZܮ �f���Q���P=�zӘ�ŤBkH#B���A����F�U5�M�Rs��4jLI�{%u�?��W���~��]L.�Ņ_������y�WS�Hc۔��M�v59*�^|�}X��"��}:��}������p��CcP������;Ȍk���6�NCH�,�#�f��ȷ�h�X���)�P��u;�j��?,TXJ
��2�"߈�e��Z��V�P��^�8�2ѷxm�@�e���m�'�z����
 ��+���E��ހ�!���qk�$%��gҾ�K�����E�����M)�H��=5}�ą�Gx���LS-)=�D?�}.^M����Q]z- ?�����ywW�RJk��\;5��ܻ&i�� �=SFo��O���Fblԕ������������@&8����#T,͵�3���F^8�ђr�����3���c	� 4k�D`���/m�/�y�Ԑ�lKД b,�d�6�!Y{7ɂ��R�F޹����Ҿf3c{'dV2嫪�ӭ�������+���zޜW��ۇAҩ�x�k�eu�(U�L��i`�>�qG��F�z��a�왳�zBE�3ig���E��e���[z�[���iz!�a����g5-�-�c.b���{}X���D�*�^��C�Y�24�U���t��#O��2���p���,�����ȹ����� 	������%a�^���m�	ڌeG�r��k�{��A��s��]P��l0�QZ=-��K��xg��>��>��z��QB��x$T��6
H����a_X�9��(��`�����Ft)�gGm�w�fV�߳I4�AW�oir�3!s�w�b�F"�Oy<I�Lv��(c;�ư�˕�`��+ع�����)c�.B,���K
��U��1|_Q�.־~��چ�5���e r�ya�w������h�<��$���}j(��
}�S.E��a�.�Sw�v����'`�Sލ��uHC�~Y���� �2�}b:앂�|�d�Y0�p=R�f��������$ą#��P�B��s��;�=��dnSN��V��;��ޜ�W=5c��<R�%�����w���s?e�EH��+L~mg�cc��Au�g1�����z㷳�S�'��죥}0���&��O�����M2�]E�N����",q�7Q�iS.��`_IS2�eh+�rQ	w^s���*�(=8M�Z=UzsC��o,t?�3"�=��8#9�mrH��:�M�]!8J���O ��5m)�KA�ٷ��XG�&��0���4���}7�U�b��;U�a���-�R�q��*՛w�.1�0�;���C���O�*
c-� ]q��&�	�A�����a�iYT����
�Xʩg%ZQIx쵺���+��	�<(�>�N{;G�)�n#S��Ltx+���>�Vqa�i�}t�zB,6{N�g�X5�[M�q�P�>�e�D�F�e�a�Q/������� C��"q|hb�0��%��ԃ�k9w4c�OHBf6;@���U�!�ji����q9���UAͤ[��.��i8 �ſC(��� R̙/���	l<���|fuW�Nple�O.žj(��_M'��� o܂�d7��% ��a��@��¿z=?�#i��Տ�	&�����L�U嘵(�dc�E�;�{��ﳨ@J� u�~�֤��B1�u���恓늱츄�%PJ�b�� ��E>X�|<]��-+�km���j�.(O	nF�yS��J���X�y)���⿠HB�E����v8	F�s`|i�>�GR��{Hʐ����k?���5���<�U��ئ�FZ��"�����7�1H&�}��F���@���S$2������c�Ϙ��>K��x�P�\e'�O5���P� ��Ǹ�~���ʾw
��� ܮ�>)������`D3�|g�&��h?�0�[�����u����B�w�|[���/E"C2�hǞ�K����*��Z��D�	��I�#�E9��T��m��M�Fp/s9R	|�7��{���}���_��/v0f@���'j/
���P0K�\v���)鍿f^���U�W|X6������o�dF�SL��Њ�b�������<k b�\Y�� דWw��d^$J&�"bPg�.ח�.O�.���D��_�u�&|��z�QA -,�hǯƏ��\��O���y�u��\�Ƃ�*zS/.v+o��2Ϧ��61+-���O���iT@���%�V����|E懿�3&i��;9Ed[8��zN�n�)�+ Ou��A/����^��ԬC�]��B�X���u��>r*�Q�j���tq±�iQڨ�T�2I��9�5R���H"�B�'�p�l�(�PÌ�i��t�(�҅��{�2'+e���uo��tn�ڏKc��G�֭���g ����?��M�4�]bD�wbI�[���P��Cr�6	'���t͟�+��0�/��,��G�Ѽ�9�4����B��?186�!�.6�,,�������[%p�H_<H@�ж���6����N���ɠ��L=�W�ƥMucw䬀C���ïT����A�N!��F�Tc��4�peq=��N�ћ֓�`O5��p4�+�"�G� �B���X�P99�v��_��h�]Ť���<��ⳡ��x������X2b�yo��6�7�?����f�5.�pf���җM�씒S�FJ]xjRy`93��?#���'�:�݃��Cӱ��g+ڗ�]��f��8`W%�O���C�ɜ�É��pP��g���h����2�y��)��TT��	k4tJ�A��J�q�j$<�ʊC�u��`}��[�i�H���`O�'S a�w��X�6<����r�y!u�h��7��)��Hߗ*�3I���݋��a� ���A)Tī���$��s�e�M���U�i^J��m^i�@9�1b]Qh2�䶙�
N�v��/��2g�EK�QJ�����k.p'�<�%v��P�zC�Vb
rz��O��b�(~���͏�BQ�p9��C���/�������q}ފ��"�6Ц���bQ9e:�,<M=S���s�s;��::w�H},��w�*/��=w<�~L�����l�2yo����e`=��̗ۢ�x�4Ls�����↓����*Mf;�$`�C'H���[2�RBA�̨����SՉ��������ҝ� �Y��m�a��ʦec�ׇ�,�k��O� �n���f�U���B3[$��[�$F.��t�H*�56��c�;u�����N^*��{V߽$��*z��I�9z���A���r�O���E�@J9Lۄ^��kVF޷��P�+�֒���O�������3�G"<���|��,�P�X�ޕ�7D�V!u�k(��H"*�Xf��JD�}#�k	�c\�9>��о�BPni|� L��c']�5D"��b���	��(y�;�ּ]sEZ��H������� B�f	Y�|�_��I��źM\�lH�DV���$j{�H	�o}��;�j]p�*��8H���sB�)�t0Bux_�U�B	7S�/��}\���%�b�'�+����̛��J��d�p+�U�C�:#��K��5�K�M�&�����%E��!b7R��=޿��8����Q1X|5��9՚���cܶS0�Q?�)�C�!�[~3��I⾆3	��V���,���CM���~B�W���Ve��܎�;�?�`x��u��~?;t�բ^,��K��+@��S�-[��5�'�`�3�Ӌ�}����E����t���]��~<���]����_D�Z8��tgu-_��N����(ϸ�{��_������J��>�q")����l�}�I7R���S�L��S�E.�&�{�d�h��("qy�F����g�| � ]���o��"M,�Ᏺ<���eQ�3�3��~��~�\��XS��=��Ԅ�rLE�D줅ژ��aqR�W�3�� �zkA�����s�`]|�N�M��G�-	(��bM������uh��ׁ�@���m�8����<��~O��d ��pJDŹ��Xӥ U��3Rd8��=(�1�Շ ���d^�1@��M$$V�&RMZ�d���^�y�xR�0�ny>����@4��~�M��"��u������B�B�i��2����p7>{_�|��n�b���e��eYx~!�;�)�5	#t���a�"�VF��a�P��,���錾�=Y��n
j���@n���qGݟ�*i@�y�V' �;��W�sH#�08�f7�Wz���Ͽw�P�:Q���R����������th\���Qx�zp(�<4x�����P���>�f�	V:���� �cٰוӫod��gSV���p8 gv����$��I�����u+��s�.���5�șN�*�R���ukOw�j�/1��xm{!�V]���2@�5��b��_��XM����C�����.N����u�u�w��
�͇�{���2�Mr���m�����@;I�RگF�� 7
���/P��EQ(a�7�{��&p/���x�9��זPnf�U�wNo1�
�����=���8x(��lT�f'-k�g��ǰ4m/U2p��#�Q�i2#�es���n�j��d�������`^k����^�.��UW4f����ǩ�5�- 8("�PF`���2Y�#m�܌�k����ƾ�GF�.�H8���t�ߖ�����������ʼ��
��_|J	2��>���
�X��oܸէ P������s}�����~h�~��Ś[W�Z4Q��u����>���f;�
VC�r��:��VC��+����M�q1��ӏ8
G���+���>c�۸�0g��L��'��쫄��v|��g'�S��+;��d��ϒ.O"��B��Z���(Y��b��j���SՕ,�Q���aĎ�-�&�O_F�֞֎���*Ff���af�EI���x%�4���:n��6�r��M�a�1�.��5S�gڢx�y@L����f.3
��w���>)��B(�W^�e����ᛋ�o���Xɘ����1�����B�j������e�QS�f"U�N+�JF�����+��7NõaRD�=���iX��ĺدl��顪R�i�D�6�/^��;��U��0%X��km���M:J�퐓�'������-��m��κ]��B�`?�=��^�e��z+l�V����i�V2n��.�Y.��߃��-�eA�ܠ?�oP���P9��d���9�����J�o�t��W����Ds2��|g�&]�^���##�[�X6Z�'�� ���q� T�Bυ�c#帮��g�-u��)��K������k���ʐ��')�	��$��5d���(B2���D�� ��p���R����x4�e��⻷�v#��`ě�+������A�:��(���&������(8���\����B��T@O����W��M^���=O�:���a�}��0,�bEd$o���(j�bOο����"���H����!  �&�߉G"�XxA]x�����k1}�
g��o:o_&�)Iؑ$y!<��W�F�z��EEَU۱�=�J{��o�KAٝ�k��������i��*�Ь
�*���c���sYfM������B�5i�=��x]�����9�>����8w��3/~GV{�$�/��?�\�a�U����J8�c(f��Y��t�l�]��E�a�V5����BF�C�(�6���ԡSv�)���I[�>_���b��Q��O�3���37�z��^3�I$%_�[_찜m����05��̮����Ac!T8S�+�bw}m_a	y�fx��N#Oed��+/A����5�9b���AQ$�`�sr�xO���X~������[�pX��3f�曠�1��l4Hvf8R�6�8޾�g�D{�a�ǃ�=���l�ӦD��r��D���I�TՋ<��Q�#NB������t;���1Lp�9:�ے�R�3��Y@G8������q�=�K�z ��Tzx���� ��]�?�Y�*�Y���N�]񅴩UV}zSS���_������и����I #�p�7�a'�/z���ʻ�%�i��(f��v�ܑ��Z{��;?+�N����1~6C�Q�F_HW#�/c���Cp�˽�`	j�Q��J�}�ۢp�!ֈA��J;*�*��6Nģ<Xeǁ�C��݂�+����B��ʖYF>�t�t�A� m]�`�1�O���7A#��tK,x��L_L��ts����z�Ty#�wG��`R����\l�P�����[�p	����I���xۂ��c܍;� \�B�.v�jҥ�R��}��n�<���l�i��A��0�n�naR�&��d��\u���wg�Qf��|)�F��B'm	<)[��)����	��6H�;�z6J�	b��Ɗ�|_�����;���tk[J�<��^�5'� }~C�꥛}�E�ON,D�[�W�tF�Ļ���Cȝ6�)-�d�`�'�+�Q$���C#%�2z 셒�~aI8�B
֜���+Q�6}��B�6�D8r&�F�xF�CrC'�YmP֯T�u	o��v�@�)[%3�g�5?�_���=ߋ�����h��c�M	�>3�H`���_����D��9��|�"�:5(�/$�߭���8�k��;dЙ��%�iC����6:E�;	�]��,1`�ĺ�(�=P�_�Uz�^9�)#m��d��{PaƼq�c��vk��V�F��U�͹8��Hi�����?���Q�1��,pŊsM����@�a�F�z��ϭ��L�oy2�xۨ��0g�_���7��ϧ��X��� ��7�(���tXp=�9����l������L�6�k�X���Ǫy��a�Z�HHDF�_Ǜ&�Fz�.�����3���.iXLCql�8)Q���n<��q��y����c��)R��f��Y�?�P/癮]KI�	p��.�7<��;�!��Q^��ɗU���UQ�����N�Z��\�mzUt��HRYC�W��#�� l�ێr�tC��;��_G���r ��q��,H���[�r8�e3}�9��H7��w�p޽� �J�ࡶ)��KҦgY�88.������C=Er�ׅF�W��օ�e�\���� ���	���Gv�mC��"vuf��<6"��w���z��9�@nDDކ���=�l��� �a��
��w'9<�`I{�|E\m�O�I���w�zT|���^2�8�����~"��W�imF!�M5z�@?�t�B��^� "�;Ā #t�Q^�!G�R=j�Ѷm����|JIS�����[�Fc�7ߒ�=d�s��mB���] ��#k*Ƶ�󽍇���쿙������~�M�"��S �lX� 6����(��z�9c�G_i��2�n;=F,��g�0P�˽D���m{�T5��4G�+�b<���'�����>OH�#%D�?p��_i�
|��x{�A��A����ұJ�짌�2�#*9���X�7F��CϮ�	��ǳ�0��M��Ŵ��5	*x��1��۴��)���"��	���UL2��z(k���c��A�^e��^C�D��,��=i�叫%�چ���<�>���Q;�A�t~�W��±b7���(�*<�h2����������2�,F���j��眔�D8ׇ 97�z���<�[zK �t�G�ٲ�-1q�����i���re��H�ݎ;s�G�Q'��56ϼ)aFD�:�˭�.��R�1��%�xK�2��{C��4o�xr�1�%�� ��G��xڝg���FW��8E�Z�0�z�ٟ�jd1Ҥ���XC�¬�R�z�1ܝ�G�=7��/t�����!����=_�2�9���G.%��Vu/td���g��yf�onb�}Pʖ3����;j
�� ��s��D�ȓ��'h���\�׼��VR��(��^���"��d�R�����z�g�t�0�4[��?���Τ>:�Wq�NՖ�{0��Ȫe�G�� 7$pM�~Z=�Mɾ�@�a�k_7m�@8��MD,BgS�>������x�n�oTx}���-��4���@��#��q> ,��$��xu0fꞾ�lS�\֨Ao��t����Zt���uf1�8���F�K��E�YO��[��ю�mO
���75H1���J:I^�w����x��V����k����H>6\��c��0�^f�
Y��{����CX�df`z��V�W5~G��u���4+2�G�p	R���ռk"F���+�8� 6V�5I�����ݘpw^UU12�	7q�%�҄��!����pl �|5`�ˀ�]b?ӗk]�*N�)(JA]%���a|�[ՑM���>�m
��m�?�Q0��{�����r/*(9u�L���6�j�"ā�U�Q{�i�=d%��$Y�lA����dS�K��I+WH䓝����oT��AR^۹�x�W-h���U��H�_YxΧo�ūy��P/;�{��#�1��ޞ��N��ݷ��a�en7�p��OxlZ]�|*�G�P�������7jO"���;�F��|$_�Z�++�L�f<�� �-Y>�9�}������6eI���
���9�"�D�A�l�Y����`�rf]�Շ������g�-"I�'�OO���#D���s��i�%���AmN԰/{�����,�}_F���0��d~,�n��`� =�n��o��
	߱i6ĕ;�F�,K��d�Ҫ\��GǼN�q��K��6�w�O=ewY�����g�������Зv6�%��BR��!��9������i�o}�dK\I�s�B���/U?��Ɠ�\�ͷ��@����2x��a��2��o`�{�#�N�@�(h��Q�t/�g���ĈT�}�-ay���PK��(Й������� ����r(��m����m_MFXWo!�g��s��z�ŀ���t)@f�1�:k�}=�%��0auQçd!��Ii��u�ۤެ��Ik����{���h(�Vd �4qsX�����w ���R��C���{c6=��DP�ddΝ���"ɮ^��Łn�#�\d�z��8]�w��H�أ=v��R)����wh��ّ1�������;���+"�,ʄ�������f\ԋ�o>�"jk:�����CG�,ɭW���~[�_6`暥�G�OG-Cv�}��P����X^�4}3�� �8��ጦ�@��*uH�ϕ���}���?�S�<2�xɕxl���g�O-~<��V�4v^��7y��d��fA��>m3�ڃ�9���Is,�ܣ��"��ᘟ�$���`���/�u��x�ӯ���FG�E� ie.���}h��~��P*%˞]b(��הq!��(��9[$�5��R�!핍�t6�z��߸��Q�q�Np=��D�d�RU�Mz���䪚����(1|���r"<��<�TC�tAc6��L۲�}���?~]~(^p�|�d|�oj��綵W6:��ծ������]�#9T��i
�A� "������4SM��_��-�QG�U�V�>��Tx���ਸ-_�ݴ��7Y�a�{��*�8�D�Q"#�|S #�~&N��l*Xabz�#ݠa
me̠6*ɀAO�n(�����6��\qh�]���W�A�K�Ս�k���;�AvqI�=Z�Jz��V	�m�SQ3�ws��9d,Y����rd� =ܥ�#6+*�p�Kd�!�'�N�Z�s���I���y�g�M�Vt�|K� |h:��j�]�Yq�46̝�v�=e�ܨ��f�����PC�%��ځ�1G6�y�y��W�V�C�"G��-[���=���t������9s�6?�|B�Ҽ��J�Cf�O��r���uc�]@�V?N�KĢ��0��|� �:"Q����a��n.��U�N��QIy��l"\�[�$�	����<�D���7�� ��ӓ������2aw��zW
$�P�rޫ/���b!tCNA�\����@��[w��[�9�������+6�#���h01e��F��<��1ngw�l�:B���:����ޝ����rZ���=�}ĉ�������	QӐ}����L6�E�.�=j�����P����}�u[F(�;n����o�@s�{��k�?f��I4҃�e���y|_���V0g|V�n�B��ѺD��s:W�wޏZ�I�HE�(��Ӡ�����)P�E�2 �S��,³���`-q�I�ƭ��/���x0�*��`"��R*.��t!��n,Ζ��
�6G�C��ŔX�>@Uހ!-��h7W
��u���(��/	�a%+[l{�2�*mUM,1�zH�{�3�3�����Lv:�5\a��)��?�JZj�'��CZ��G9��+���ɴ��H��� nX�r�5ӯ�7� �Ō��k,T4SU���C�͂��D��L���/��=���AeJ>\9��Rܽk�v�~���X�^[1�������G�h8��|F �<��QdNQ+ؒ��ZS��6��R�;��	����Q�.Ml�8�N��j�� �҄!�s ��!�o�	��)�bLL������p���`�/����o���h;'D�eK4�jE��ȿzՇ���+���wܠ6_0��Z@JK�o9?�
�!"c�rM�v^����h���3B��qq{]��9矮�&���h�f0�~�? ����"L�;�]�U��7�svC5ݜh���4��V��i�]C�;꼔�]��}i�<G,��ڣ����[@��u�i�J���׻Jsڰt{��g�b�?���	w`)���g�16�l�x�[��v�Ml)`¤*t�S�������}�ᤝ8���:׃�KŦO[t���Cx�����!�n2z�3�¡����N,2*q8�o�	�_��g���*XyfS��6���D8���Z�:rZ�m��#��u���d������+1~ц��z|��%���_��)�mO,!U������b�gŴ
�%�<�����[Y�� k�飊�m��2��4hj�8|��[û��A�(ߵwD
��!딄%-�vʣd�@�3�&�$��o{{}B{R�o�ђ�7��_�����7[=ݪcj����L�����Ѭ��"Pp{��&J��`����X������C���2{�j1���Z���S{~
���T��O����~{H�&�\�$z#���/i��%���w��J�ʮ�ue|x�R�l�!��P/��Ɩ`��o��"�n2wJ�G�|�n�(Ɋ���p�;�x�1�cQ��n*���yy�����ő���-��_\�ڿ���2x�cL0�<=��R�Ip�Ѭ�A<Q����Ϟ͔s^ ���Tq��B۝~�Nǩ|�A��ilm�C��|i��)gg�*�!�El�賮;�΁�&΁��]2�}W�A�I�9c�#�/�q�V�����|�(�~V��+��cHY����[�m*>3��?~�+ս�D�:��^�}����Y�6���&�� S�Za��	%�'v��@E�ʮ0�Σ��|�n���y8��e��-R��v���!]���&aJ�!Y`d`�}d���S������J�Lڠ�zF���RJ@����:{��	���ٕ�����ԅX=��wğO"Z��CV;��