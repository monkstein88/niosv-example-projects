��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���~�`���sB�G����f��F�Cx�2��ܹU�`@?���ٚ���y5T��
�)���2�*�O;�e2"�_����q�2�x�����،ȱ<�F��e���@y��'o�D�w��X���oFU����c�$c���bM���?@�̯��|nY��T�;t�b��T"ȴ�Vw�D�W{�c8e��%�
%b��0(���'J�6d�����d���cq���y	�Cv5��X�m��X�R7��eJ�g��Ȱ����Μ��9�G7(݈�z_U��+����#��Z�hi�R5���a�&&�w��J�=�?�Z���o���zW�G0t���t�����dC^H��������ĂC2�^�6.�<$��Lqe%I����MC��'ΛXGF�ĳ��7���\��%w��֛�K��(?�;�>P,ttuB��d�o�1(�U�4���KW�[�"��sI��Y/w�S>��j_� �����@yLB���g�.Z��g煿O���I&oF�M��p����βa��ԯF��o���q�WtI�4�!�C:f&��a��6�RE���8L�:�J����\F�>רxS��e�n��ԟ����=eL~� ����k5ȭ���(4�⢠Co�~���Y��mp�;O��BX�N�U>$�����-E��>�&�O�����w5�@1
{svl��
�Y!�p�x�r0���a�����!2�2�.��R�}�9�hr8���".}����W�9�U���ޱR��)�m9��S�=7=9�A��گ���퇱�ر�c�d&m߫c��A�XGQU$i�5�Jv���O���+�����.���Ce�ߤI���[�9�����,�Al�6w��SV�6軫��U��rr}"*��ZA>y)�����$S/a@��p��x]=��/jF���du`��#�}mt"!�[�̗�Y0���2+Dq���	V���)���ձ_M��%��c��[mv����k⤬3���i���l�G�Ti�K���7b���|p*�@�	(�,tI0�Ă���l�	��� �*.�f���7ɑ�ׁ!H�ߞ��޾�E��_S�OA�5\&��JA��1�Q���}ϋWtX'��I��m�U�8��$.U �'ٷbq��%d���Ew���;V�1Fyx����*4d;��Oi�f�y��D��C��ZW?��.�,Ҩ���R"�/��X\�|��y$�	�1�pL�uĝ9��w����o�
�8��e-��rl`��!��h��fN8���4t�2!�'�]�c��s��Д9�/W��a=����?�p��*�D�pŬVea!4��^���rE~��!�X���Xuh��뜍+�V�̘Ui
����n%�~�5��\"a�,�������Z;���#�ppl����Qg��%"Hg�z�#�02�)UwG=EकF`�A�*�!�	](!e�!���ÔC4耜��[}�@H<��IWuosӱ�G�z�CDk^�����R�Y�`��Y��4[��NJ�ݒ�Θj��[?�}��-�_"��V�3:miq8��NO{S5����[�g�c�yD��U�K�v�@��X�D���XF�M/;��D��,�� dN�s�S85��VC�u���8ӯ�I�B��@��R�	Ń�&��-[��S ���pVX`p�2#�S_W�ɰ��Z�X�3xdV���������	/^�/Wj?s�a�M��1�[�\�(���bA"�P�VfB��;��\��1�����z����02-e��+o�}��{g�h�A��{b���Yv̽]����T�k��pF�����績ۥ��#m\!�f��b���)���9RD�^9���o�e1Wy�A�������/���y&;Wya�
}{AS[$ѻ�2/c��{��P^$m���p�ٟP<�?����&,Mn�����dy�n#���S���.�e��R��\�{��*�I׾�pw��* �6�fF\�aW`���ѫ��Oq�/�=�K��R(�廀��Z>ksho���1*�jD7 ��e�o?4`X�ci>7>����� <q[]!\ƕ���Zl%�E���B��@���X�`�&c��$�/�k�ݢPS�F��9|� d�-��%L���Y�XYrrAM
F��R͙%hF�S�)U����G|��ڑ1j*���%AMIkD5�xU�щ-Aʚ��iP]U�Q�,��V^FV��/�΋�ױ�U��e
zm�y�V��l���t�/��Ҩ��F|��2h���D���t�g�ϖ7����#Ƕu�K �e�c�@�y�����Ŋ�vAj��&gv���w���G d(`m��ae��8V�'�T�ۗ�~xm�/���x�$�F���a2��<���T\�HȀ�I�;UD�_#�i+����D!�):��C�U���Ɗ�hi�ҍť��7!���f�D�)=3��晏%���h�^u99,��>�(߳��pz���{�&�e�e���t��51*��-fI��f\�2~�%sb Q�[�6�'e�7_}ś����:�һ�r��5���/�1��mb�ߛ;װ-v�N�p������X���Go��j|�"����#���E��v^Z��E�ݪK>4���\�{���UA� ٱ��:�$��w�'�a�&�%ZP��5bASdֿ�$�r�ӕ���<2sDo�V��/���~T���0�?�IX�g�|�B4Xpj��N>�c�|��H�
a*0	�{�h5~;̼Z|c�]���� R$���e��'sy��\gm�ci%]DG�F�/�g!tֆk'�5Y�L&��⠨ж'8i>�;�ވ�j���vA�%�5�g��Y���1�mIx;*��"�bX�y ���C!���ܔ�KMs���o���8�N{�ੴG8+`QY
e��۫Cg���т®,f�Pv9Aa7�TO
�).�3���Q�������N�:�h��t���=�5����S�"Z���fJ�~��Ĝ ����&����@��3�{_i�dV7�|�2q�VS��)�{*�w�
�;���Q���ˮ�8:�}T n�Ъ�a|�3~��(���V>�g6�D}�й}�[U��_'�y�B�C��Ph�GK�c�2�egRe�M�h|� ���K+��;�$�}�TV�ĉ�����Н����p@X�h���O}qr��8"���i9i��
D�>���%A�W��i��6�W�h7�B�Y_�]�F�ԣ�f1��ɥ�m�|*�$Uots�8>��z����p͔_���~N���/���{�1�����Cٜ<[�������	� kf�H�#jFO�A�oy�S-��g��Y�=�F*�w��<Ʊ�"'���1g䥯Z���_ߔ�m�"�G@}Է�|�3����y�����������|��v{�d6\�$ąB73��z;�/a��e�ԋ�I*���
��u��Z�<���D�JϚ}��dDp��F������>���r�,#�ڱ�f����"�a)��7��g*X%��C\�?hցC�SS��߂E6�w-I;��Ha����Y��צ@ֺ�����Eh��R\��$���Vk%MYfa�+�e�@?���9�uk���B��z������9`����ӟ0��6��W�4A�h���2�tt��h�*+ ���b��z�0fu$@8�ه�|uǵ��h��6���H��(G�~�U�X�B�/��-�r&�Y����)��y�z�6�T牽?���k@���� �Us�w�Y�z��?Ǒ��(uЏ��ؐQ�[,3��1�E1
�)��q��Z���r9�خ�mO�kO؛¤xDw����UVΛ�~^�[�efrS-P�~����E�D���?qX0u9�YPC�4~�Sf$�Q��'���)r���N�%�~�&�Z�ˤʖm���:�P�����#1�1�G���FwZ�$!!�Vd�J:��jV'dcBQ��l�K*s��B�S5^g9���ñ�~ª�x��5�4:����l<�quD�=����i{�'�Qp��n)�E��J�Sݙ@}:j���Qu���\F�C���_���_�S7jq`9�"������a��{t>Q��ĕ�%gF�&TQn[���D��c�=�<��^�5;NVB-?Yn�rvJ�]b�a�B���1[T��]�R��L��K�#"�QgbtÉN�R �*y��Vо��i�nz���s��J��h�mZ�A��W��+0��|  ��O 	 I����9C��t'L"	�.J�q�~��V��@:������
%RN�ن����?O�����XG����/��ڀ�ΟL�4S��A�~F�9.
4�W����rz_�?X#j@�)Ã�&+�~@u_q����Sפ� t�y��|�b�YG�\5�.�"83�΄̨?v�.0x��S)�8�)D�<�<���q���7-~�sz������g�|"�#�S����˯���%AW�	�L;��5��=�J�i��Y��݈��x�hcZ|�q�&
NA�_8���}s��܍�ԁ����f���ܗ�3bEӑ�,�����1������r��3�n�M���p(rhU#��AH�qyH���V|Ï��y����"pŰ�"Zp�I@����P ;at=������{��I��º�5rH��$|�JX�_%s-X;��#�a�+'��(
�i�����En�E�¾~��"r ��ɰb%���3S/'Lz���etฬ��Ҿ/>�~>�Bɧ�4��|V�v*�ג�����$~�L���������ƔΠE�;��bj�G|�6�0�X�n7�\+ۉ�d܆�68�K�A�e�^
xl~��bV��uN�r2�"2AS�11�H-r��^ִ�%��Y�^EtD�.���LT?�Cd�2�����8B⇒�����~�O[��sC�C�Rv�4|[Uæ��|Y=r��A#�h�\��6�	��U��_��{4G�Zt���GI�bo�L
�ou@���#v2NbR�mv��{/�����$i���p��svm^r����c_��к����Q$��H��f/�q�?4e�Y`�<���m��7��C?��{��bǥ������;� �@�ƗH@�U�D��ߟ�d�����n��"�*���]��k�A�)E��u�DQ��;`U)0�(i�BC_�俽�' \�X��56���5�<s��mih���� P�Ȳy�ߠaw�%�\l�����~��rU��z�C��d��'_��>F����3�l�(�z*���dҹivr.svtߵ�i9\�3�y��i�k��qu�����_e���A:w#	",n��ޟ��rȇw9(���d�R��a48��l'uo����
`�A%��ao�:�
���O�҆yQ�4p��.�|39mQ��Q�ӢY۠P��¯�@D��j�N��#Ig��_xgK�T�3��g��Dk���t��STgdpR�b�Z���[R�U��x?Zv%��e�2p�B�M2�*�I�?�jQ<��n�y	D�7�c��U��Lsc��`������@�ϴ��7k�څ�q�Cbƍ���~&��_@"|�������vg9�����.1"0�����w�h��ogY�=��9�� ��^p^?r�>v��"�b�~�U�#��9�Z�w |@1xw:A��"_`7Lb�x�������;��9T(!�`�U��4��X#��Q-�X2m?�����1�=�['gR��%��Fb����SRvi3�-J+�,U�Q�ƾ�ؿs��&Z����;�W�*��j9�(i��W��E��do���V1"� ��v��� 6������F%�|x1��B	��W>�����p��[|���L
O�;�rá�g�+�A��T��i��j�t��|ռ��@����?�k{����Y�F%b��$�y�W �O.8���k��w���}�g������TxP$f~˾:{u��?I�� ����Q�#�>tF�`2;��U% �w�A)Wx���.���KF4�ⲟL�b]ƈ�W ������?$�3v���r|7i��^H����'�3��9<�R���n�bе-��i�D/�(�����@6}���KRo�%]Cdʅ���C�����G^�G$R5x�>�SɘuK�%��
?Um��nw��1��K3�0Tb��P��@�ϛkw y�����,ް�m	�a���k��*.+��8���
�6�5m/��脌��_����L���`%.Н�S]?ϼ�ȋwC[�o&\���y;d���2�a�������7� �y����B��fYe�XCZ)%3W����Q$����&�Om_+P�	��7��&B���6~�H�?Y& (E1��$�>p-���:�Ծ���Y�'�������MENC�7��4iL?��q�"�L?��]��H��ͅ�@�5f��(�,�g�&��2�K\É�V���?ؚ���Hd9��ݩB�9���hl,�F)	���BXer.L'���e�q5�x|U���j��qV�ZBU%>|�Ds+P���f��z�`5�