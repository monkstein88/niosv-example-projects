��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a���?�;��ȎɌ�K�-B���b��Ƚ�/'��{��> ��	^FV�X�;^iQ;
x��}3�X�R��/�b#�x��*�"xH���M���'NX�䕇�,�{��m�D�\�%ߥ�$�Lo�:htuR��$E$�! ,��gm�:6F��1%JC�� ���uwJH�I�"w�e����o}H�Qʿ@'�1��k�l�ÊF
�G1����4�c̓�u�c�E	�Ԙp�r�|�a���w�7j�n
�n	�	������b�Q�����x����!09�\.K�ݩ��Ǳ�.U��9{��b@ʠ��A{Y�� *�usMZM��0q��:mޢAЯ�)�+��I���5�=6���Y�S�e|Zǧ/��:�!&W�wg�� Y�}�$�[�	�b�~��Q�zZ�pOJ�B��ݳ�(r��PHj��@�y����-X	�v70��Y&�8e���ݐ�`�'�[, �������,��K@D/��8!�����@j�6��+ţ��yp�����qh���+�J^�J*j�X���d+�j�'F��l�5[z�!����dnAe�����%QCS �L40k��據 ���$�9aȣ��nw���yY��oܬI6�*��a�����8-��mqo�x�)�5)��Z}C�h�D.]�Ptr+w7���ь�R�$����G�׷�Lpe:�kS�h¤)� VR�(�O��)l1�b���⍙#=)q��Wz��˿���)���d��
�h�S(T����;/?���G��/ɗ��+nW����3��	�g,2o��Q�}m<ڡ1��nz�ǻ1�ڴy��D���Ծ�"�(�f�VY�s ڍ�yY�pՇ��d4�r��\2P�b!hk��4�N� �ڏcQy�]�M����� ��Emy�lE��>,作a��b�Ch��Ō8uϹ�#������2�L_jU\	�/n!B◻Mt��%��K� �8兂++�d6��U��i�Q`",Y|r���U���V����l�_׭�3�f~�l�_U�x��0�F���%�����?��v�G�,	:��!ܧ�Y�a�}2�168�;05���΢��8�7y�e!����s����*���T�� y�\��<��.���4�1O��z�6�m��N�<�W�����зvx"�z�2GVTs0�T�6I��{�6c�lXN�A����w�a�\Gd+�)yH��R��ee?�tW����yAC�?6�ek�4��~��_oG�CG�Γ����6���DA������
�N�q��R�s#n�*'6���c� )Mż�:!L��ѡ$;�J �\V�ٰ��r��!Fi��A_H,�O$�_�S��q�*�Q�t��S�y��wb^s4&��~	� ���^W)��u%��Rq\u�Y�*$5/M�	�'�e�)��дO��L3�.��Uj�=�:}>FÜ���1��Fy���� �&Um笙JԶ��4�0*�0�d��X�B :�+z'����hj��a<�� `�"����*��U�����}<�5�]s`m1[�vNw!c�h�X`�Nr��'r��?�~Ɋ4��dx���Xv�Z�U�%wAaa�|'���z�"�tT�NG9 B+�d^�A:3j���u�뢋�cp����W	���yH���5�p��И�ܗ���<�l��jƔ����mb�@�K��]8��z�dE�C�[5�l"������	�7�ކ8:�F��io(��s`cr��<T�hʠR�2ƙ�e�vM!l�,�JS�^�?hk��e�ǻ�w���:ON 9x6W�s [C,au&��jE�0W3V:�O�Dl6���b!��%q�I}.ص�cJ������`oLal�ʉ',2��Ѝ�\�؆]��T��>��w���W	������ �Fb�3�)��PU��wbı���n�������<6R}_�����e"#/�芐A��#ʱ�
��B�In&h�~R�;z	e��!����o�)~y����TFwh�6f��G�={�rUP.����\
m0���y��nn�:fa���(+�>\%0��H���g�E%ej��!Y#�]����q�L��ׁ=e��nPӔm���mM���,7�qro�K0Մ�äk��Ն��o���H2d�������*㒎)9y���m�,@ V��R돠�.�-�*,������<}���a�R�<���{�(t�2�r�d�?E��\��o�t��[�y���<Q��M\��I%nf#}`s�  ~�(ټJրhJ�k�y�x��ֲ$���N�sB �ՊB�!.0�>�bG�;S���t��J�;:v�o�M���W�z��i�Yį�f��,�[0��ba�Y��-�Dܿ���:��poE^��=��C�Ci�@?&�������Ǔj��$\'5��3����7=���ɏ�w�jt���gJ�зiW�'��d�,�5�����9Ӥ'����}��5��v����x#ͫk)����ݯ>�V�N��)�d�Y/tk�Y��߄`2�p��r;�"Z�5�}��hv)i�X��owa��{�w�}���{k�I��h(����#ͅ��f	�\�@\����_qg�ȧq=��Ɲ~R$��pu h��c�( �R��X+�v�ޤ��vW��\z�zd�9���ֹ�����p��V!��kR5"�T�3JKiS9�8��fJ�і�
��h�c�K�ȸ�ލ|�+�oS���˥���u��.�̞�a�C^����������D)Qe�H�hbpE7�B�D�>4l�_W$��G��Ӻ��b�d·-P�{C@��B��!�p��-(==wŚ?R�78B�2ޛ����A��n���6�����0߈��;qѮ.G����4='S�P��8r�l��(��8.���7g6c� �C�'ua��R��PI	�� ��J�w�EwMxˋ=��e^�bឬ�n_����h���Y���3F6���")Ɠ�u/6�E2:���l�OI��2>&�),Z9�"��Xy��^�j�\�������e�4�+f<%DG�F`ަ'��yш�Nҟ6J���'�4�U��N��ŝ-fbl�`�n� ����=��<�\Vn�r+B��u�h�`J��b��e�U�gC���qPX%��*���jC�H�ϫ)KCıf��17�C,jP��-[:8���S�HxI�՝�C���2B�s�Z�F���(>���l���@�V�~e��[`���oO&����n���f�?� �г �}؍opUw�wm�G	F�D<�z���yȅ�|�Z��j|J|�X_�BQ`����I�yĬu�a-ϣ���>_����/{1*���ƥ����26B�`t��LYGgT��̒.@1`�2�l��;7~��F��~f�I��4���C52Za��(ʓ,�rxl[�SY��p��5~����6¨����v|S�o�~s�Bv�>~��,_u�[��7Ѻt'��,8S=ER�s��~� �z���&W0����l��AG��8���M��/�@����/��>��m�W����a!��|�y٫4����g��?M��p����WJ�~��t1���E�}�y��M�a�'�\	�-j�ԟ�XS}폛���	#M��mqbȘ�dmui�&�r��qi;Ӳ���|�:M�e�UjT��_S�Ŕ��[�?0�(u���I�;Bx'XtQu�v�>my.�
Z�XkP�e�����y+�f�A�Ns�C\���o��I��Oy �(G�����ƛ/�,��щq����T�0����L�� �bo��C���߹*��$�dM���N{y����n�"���֠���������,eJ�R�)�>��)�����H�\�
UoV �6#S{l���u�h_M�%Q�Jz�h�Or`OcV�4��cg+Ց� j��K�؈N~��A*D�\�25_X��%�M���_$�[��l3���,�+��XV�|��\�T91m�G��(�޻s��	`Ō�4�N?�&B�X�_�{7���*�%兵�m˴���cdo�4�C�[~�I�I�Zv:MQ)g�
k�&$�TRX$��"������b�a�x����&\1�7]��	���[�;��z�_j����7�^������(4.K�z�ɗ��&w�.�&�]�Xf1*����a �H��;�c��/'��Ҥ�뜎�;��-�
��9M�.��5��N%�R,8i����6A���	Yș2�S��{�٤'�M�jXݻ��t��k��Dd6�.>�?�U)��~���w�����c������=�@$:udeH�:���ѭu�(Q̛&���c�b�);��M�F�is��\`
} Ҹ�{(���rD�NLe��1�kK�Yv׎��J�������� [��B	!~���g�xʱ�H�!�HH�������>0�e��bq�{+�x7;H��q5���@B���ѡ����B��`�@�JI��(q�� ��w��|�EXos�����t1�x����������7��;2Ɏ��Nd��߬-p�;�cX᭎����M5�=��x2/C���4�ZϻA�ӂ�]���鱅��9u���u�ݳe��r��Y�AD[,�)��F��զ3�~������3���و�U���	+���i6%�K6s���41V)�b4ӯ�c���h9|6t�l������U6�S|���}�P�-���9�]Vo��iH���
�d~k�8�ᖧʎ#)����*	�陕|c���1��פ���Lm�$!�8��1N��/�1"�/��g�%"V
�[�<W0����(D��c�*��E7�ķݾ���
P
��m�Z�K��3��8�r�㓠��&��ܬ���/k�4B�B��`��^���)Y��3"����+v�8s%�44�r���T�M�j�Q`�HH�˿D�=V`0-��Y_zT޴Яh�LGpdd8���	Sh¦ojL�q�n��*�F�fǻ��8�Z'M��������r!m�&�%������
Qa���1�E׃���k�R�����?��w�V�DH�pM�GUIz���n`z�ܨ��~)sA�s4�"̛�!��m���%F����1�!�Eųs�g�來���z�jK=U]C����Q+!�-���}��� ��E}��6-�^�?�\�
	'�4�Un�"����g��K�b�%@hˡ�� ���4�ο�Q������d/3C����cw)�D��P�}��q,_��N�d�<��(���~��B�{���5�Qҫnm2�%�Jvw
�
�>��4�8mRk!���;����:���aǤ'�p4����5$"���g�$D��x(�S櫆=
j���-�vKa��AK�Ȝ�Rd)(�� �RX7<�5��hu��|��6��Y���^��pntmT�l9ߣ�-F%}�E�Y��>7�o�i�/3�����mV��(�q���9B�
� ��[�dG�?_�2Ke�6��g*�� N��XIq�5
��l���O�I�e�N#0��ʠ����|Lgα�$ 	
+����M��R���W����
�_��W��I�$@f&/tX�(��`.[��6$�2v
�r�s�Oa�3P��}=�Ӌ}7��Ҍ�_��[r��t�q�~�*��k��⾺7#,�<��i�?QןO�f���\��XTh
�"35{���NW>Sv�E����2tޢm��6g�+�f���;~�߱Vb�i�z�l'{v��������)>��4��YJ���hFE��H
�Z��tR��m-^�Ex�
[��[$�?/�է�fc�L=�5[n�^���r�a����~�Ir�^��m��L�4�d+�	���@ߧ�*�.W��O�j������:��)]\z�a���T�4J�K~�Gx>b�,��+�E�)}�S����[_a�,~�v�t}��L��o�{��������q.~�'��[�%���R)��|�_�o�if %�O�;�$|;7Z���xXp��$�.��J��lj���dQ�<^OW���[iAi�F^��j�<+NO�A��l��Q7)���2~EhD�1i}M�n)��s�mJ�{��Ii�]v ��DO�}:e�,T��NrX��:Q�2��[���DWQ�VK5g�������Z�\�_���<�#��"w�POɯ?z*�1DF����'^Xi��$�6��D�L�2��hЅްB�	/HS�(�p5^�`Yj��~�Y�:h�,GOq!�vĢk%�~�|ix�X��,�x^���J�ĸ�kc�ڃw�G�w���Z���PsaT
�U����0�U�lÜ�'������@U��E�$��y3�ږ������^�{�>���h��6zG��39�
�wL]�ܶ�FQ˟ͽ.,���(�N�#;��	)��b^�h*�����7��\8�WvY���ۉ,��
��UI��s��~��#6f�*��1yO�pܪ��d�n�_X��ԦTk�}!;O �/�cyo��|�"-Fqˌ�\�De���5��CW�͂�KӦ�y���W)���L���$��6�z��n�R&����
�<a�(CK��GzA,��X	y��Ƭ�$��e�R"T��eOE��D�Rvh�謇�^�d����a�y�|�!IQ��m�������pU��}
f�h8'�A'*�����|�-I@'W�K�vv�;4�E��*�ͷg��i/"�l�����k�UI���e���|���3�g]A���-���ԩ}^lh)�?^EK�[M$��oF7�C�v1E�WÒ�]����@MC)3�`>�ٓ��a�A*�g�}I�;k����J��(��ZX}<��+y�{]�׌�­����]	���K�<�k�vb�3**rs��&]dY�6��d�=B
��,�pأ�a�4���̟9"�	]X�L��N�bMʵ](����~W��;���wXc�� JY*h�m��eqGo�7UK��W4T�aGR�����ު	AS���]>>)!�<�We�m�~������^4�r%y�(�(��Q'S�B0�����p���j��ҹG��C0���G�Z�&������x����yn��:)L�p��s~λ��k=;��*�
/�%�!��o�J��r��s���GP+5��sj�:dl���&�6�@L��;�=��K�E�Z���J�?��a��ݨ�?�2���h���d�Uw��V�=�R�n\K.w�
��ڦ�r{�R߶�'���!�c� �\��h Y.�b;��&8�`�8
�>m��J�wzҒ�R2Q�=㊍��"�<�Ȯ�h����m����%A�d@�r��kI��	�]���ɫn�����{f��d���{��,�S�?[��ŉV���� �nT����+�:����_�,(#?��`0�昈!]T��e�
N�Ɗ���ʄ�
�~b��%&F�T����`b�"yP��6� ��_ʂ1R�v��b�\�Ӊtl���o9�?�"��/��Y%ޱ+d8�?*F���GǇ<i��͛�Z�N� }K����p�5+<ڔ�%�K6��抧�O>�JNU5�i�D�3�)>&��k���_����c����w�S�9��o����)� ����}ݭ��]� �e���M�y�����{5��8e}eq�1>��8���W|��h�7f;�W�E����LRG�A���~}���G֢���<&�D҃I$�E���l�J�s���sV׍�T>&�@����&��I�p�.Ӭ�ib|���_g�V�jb�܉� - j5 ms�&'Ո�L����"7�`�,�R�	^v���K3�߿v	��Ca;&Js�BpS0�>1^S?��.B��� �}��X���%:�! K�p��|��#���Bw睬�5�U��\a�D��AU;���{Z����/����]�g����ZK�cgO����=b�P_h���P��g�ܸ�T�g�6C�}�{.�ǾrZhtc��ʬH�~	������4�"3*z�eѓݟ��&�7>7��D�z-�$��kk�b~���� �4����+D*���iv$-"��b�y��p=�����H>3�It)��'��	�X&"��&�UlR�T	(�l셦��8c�S��
��� ��ϡ=jڹh�e�q�)���F˱�1)v�����>џ���βl�z]���R�.�zi#1�<�4�ؼ{�,����*��@��+�T���~�k����@�a�bb��^��t@�<|������Y�X����a�L
y.�F�c(�-cKS��sy�0C\�V��#��q2�m�+.�6pz�/�����7��� ^��zit�F(��V��m���<�	Vvn>����8�Q=� �l��Tl��Gx%���/��m����LآMϗ����T4����	��M���"�A�{�e���l<�:po��=��㈶�K��R��T  V��7�oǙF�v��Х�k2c����zE�ŝ� �U�8�T.)��F͠%�~4�Q)u�5%�A?]���2��. -��(z�Y=E���k����ϧ�߉K�DE�?u�o1iD` ���.j��?��z���76D�|m�b�!l�Ȝ�
���g��Y�՚p�Z^A��Ţ�YQC?��s�,ƾ�[����k�Q JQ�O�]��l1��szw����B�}�dg��Ê,�����ݧ�n]S���ʹ1WA�F�(����[�l�L+R߳��X!@W�R)M[z