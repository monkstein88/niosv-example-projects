// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
NjzbYHFPG9iBDD4tnUZcxd+AUlx8cgrHpZ2bNvwA3nzWgiwoyn16r6Hj4FC/XoIqOEbZw9bYDzrf
//3e5T0EcvEAjuf9/Tlp3V83rwg2GOV0KWocl9z0Rt2ybp3q3wRilucTUd3WAvCzqkF4pXrA+nO4
UyTLHkkaPKervlLAzhQWloksIicrIu40OgJDsGi2R9LpCNbaQDNHdBwsBlos+6qRw9NUv7ZnBrmW
nYy3ib70jyE3w6ArpNsqdapo9DGD8eYf9dNroaeZZkIppWLSex1bvPGlsr0Gg2g1RyFpmzDQNt1b
hMXjYd26ABaeIldgY509funHHPEe4gUNgzDnLQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6288)
C2gJZ1VOgMlk/orf7/nSaO2TP5jIBX3V6XoZ2V8Jalgl0/C1+A2Iu9wjJhmH26PtYiK5N1l6jnxn
aWNPULsMJq9lhYilRs0BeLS5dZTkpfPGZyal7QOwciuN0zpD2YTByl7In/bUiPpCCy9KFd3OaL7D
Eb2xHBi5S/1IJJLKoMIv5MxcbEcoYpWz0yaIIX+VKqov6eC2auurF1DTEMhtaJ0vBd8ZFkDgIdyM
Biod6eG//LKSpK09Tj0UYWM1Dj6G3egWCCe3+onTLonYLRagVQQ9pKK/fu8p3Eyj21mtR/Fv6MMN
ai7g0WvM2DsHpI8mC1rdokD2326rCIX6MIlr3cSZhYMJhcjKiYXfMmXShRcbCr1Tdyoz5bxRFe1U
heSyJhWU/deTTfulhKxFMMiOEodjC7zkjtddJkpS2udMX/H1Tj+wwvNGbqmMKzbZznfEmXjBSde/
IkNh3mDmwEEieZMh+1Sqy2Vp1XHmbewvoz79CF8agZQxIYbmDG7cprDahHQD6T63PMYD1Q8oJm/m
iheJPrSPj8IAB7uVOh6Q3expLDe6fn16v+Ef1HRLO2rlmWm8uIFGjFu3sAHb4pYHFr4aaER5jUu5
JPog8tnPfsSyzJ0nLsz8MAdYSOaZomySADLvLqxNTtr/a8V5Ab3k9/7OHJnSEcAO67iu8Cwm7L3P
CjZb5iUW88XJjV1WEJcjIyQyu/rqxJJwOriM5Vf3MaRi3DiRz3gMc6BgDyGjtv5gkXPbjMUMj4r9
mx59H0N01GYTlPNnAbc8m0JIMGCjEVNFX6seZlofuT4Gz9xszasKG6DG4NfvqmZE6pBqa56evkWr
34udoEvlDBKF1D1S9cyhg57aQldT7snuy4KjxoErIIcaUELVUWoq+D2QRskEeshg6yX/S5i30KW3
mQmjNW2gxxvPiIkySFzLK/z+RRJ2NSyEOB6MLsfE5h6NaiOMmgOMsKNFEn+p11HFzXg7XqVgjpcD
CVuozCS3g99fedjQuafKRSzmUmK4Kkw/FrIkKF33t/AausdFVsw4wQrAazyqDpsvF7+q8Mcu1zEy
KkyFmuJJVW2u3N0WJTNTtxi+TD0ruU5x9KQj2wJ/Cx0wWCkEhiXYsb0+BNJZ+f2kqRiIr13wwKQz
0ZplV6njZUCgpMz13IZZ1L6QVgsNYTeCqYnItIrTnd9g0nHDZG1v0tqAs8Y6OMfnFEP5In8Ee8DR
imjJsG8zIXrz07pfFWdMa+eAuN96Yivz5YSOcrvS+rFCLfYg3pNOC4ZXrvSNlMIDLto28AAfHMRl
mmUV7gXI3VZztYmSj/Y7Dq3pzOzZo3JGYn47xmP5OQGbr9qc6LqrDcD+S9/DHoIgqyQlCI5dAwZg
7vqh/90R+AaFK6xE5i6UXOaARpaB9ikcsEpVkJ63Fj/Ai6piWX7SPeO4rS9x/U7VoKg1rdu2HHU1
PMBa3KzTCTTU2ltIErHGYtm3BzaHpZV2Woh2gGSqPdL3TivN8+1k67dPdKbb38DSQVP+k24TCQJp
l7UG6agpT5HgSRASOnAbU879l/w2gY4LwNxWuUyJNDZRH/t1k7C+uOQ0g7KURWjMsZxq5UwXIqtk
XMzuaXVNNtF5q7SDiJIHA/fuZOVxSJdVT2rErIvP8BAJhBJvBmSH5VdpSiLTQW/7K59jVl0TJNy1
tMdrshTf+lp60N2fLehkcGodOD+Pi72PDnsOgwZOcgzrp9J97czdJCjIFUUJIYY0guwhI/x6eNPa
Mhlqe0jhTw11j4QfPqGtBKjQ7CCI9WXzxkq0B/TMzpspCqvTcSKl6I/9Iamy0PzNj6W/Fav21Okb
evj6yFvY4o0cSHzAHO19yISFTum6oyrKrJB99E9xTCkamh3YrMzIe7PnSqzUiSpUspN5gQiUHN3J
LuwRufzTaygf42Bj2tyU3t8sfcaCE51CByESeNmdixNJKj4s49oeHC6imVrd95iuQDiiYMXmqspT
wmhUDDJW7NB3ZFhfAmWT1z6lronJ3JZuzeulPSAi9yfcr8tu6jsIpE4a2wjLtSkTXdPzpw0hvOb7
pMHOWILhHzOfVcH9auWrOdc4yqI20ktOFtY2KfU9dagtjuC+YNlrfiLGsjnCk+lDYBKvz9wye9mS
rlMG027WXbU5TWAu/sV9qer/lEMs0nkMtwr5JnbzPacVCczN7h/U1Ke90kqjMBlXsHkuJC/GbSON
Z1NvMPASrBurar3DV6VAsf2FALE0eRw9WXg2M1FyGi7d0stKtmOICxxCLidTt99GaelJ4e8yrc5F
FlgPxF7ZTvgPII1fbW0GosGCkB+G0z4oQ7lI258Q1skb1QbIP8nM448VZ+AtkdmboFciwQDhZVuP
AzK4bDp5OYRRVABA48ocg9O0hEOtattwOJqMaCWSLcSm9UTo+64kbTJ6boy8bjoZsP7NqmCJkjZp
9588NXd3y1NL9eJa8+z/Q5mp3yUARsQReTf6FfXr0IpCK8kRwtWGpP8vd25AKgVndvk7cgIzODt/
OsYMv1hsoQQT4SYqz/psVbq9Ji+VrsrKrZGMhQRyGosXt/DhEbQi7OSzt1M+axad4qZ2oEOlm4Y/
W/CC5N56iGNHZXaPb+6YIY9QMLxH+PPfC8SZ3am+B/cLKLw8d919Nyiy75sJkZS15D33fY0AuBXG
Y1XNZJu4pGBsNCXjH0HYGONMe6HGF3dzdOxS+4je8QYEi62zWbKbUDmXT6msymPpkA9sAsXbknJM
NC1zu6x/tjC6EnrXlMBNvWvEw2uPgWikx7KfdmRyOiXPOP+tnPf7qx+NyXNqdy8oZ2wM7H1h4Ug7
QqlgXg0BfUHCMuI5mSkx2kghOU0XeynNgCw9E3HhkYFGSGKc/ZJOYfM6kx3je0zad8UrLHFbr/OE
bu/qS6Ltagl/eHFImCbwq/PSOSyXn02SHpFciq9sEePmeZzfRVF8PXYaIvyqVrNjP6wEUtXZuH6Y
tD2ef8lTs15gwSXn0wOonY4/vO8xSBW/t3jC9OVk+tEcHMAPjY8XsgutoW7Ic+NdU7RF+KOhLy3e
0wEyIsaPKT0+wdFOv1zvx+HQWFgXYl4q3BXkZadziy3uBMvj5YshNQ8n0XGbDPSIcMVFfi8BOlLy
JW4KVWHDuQ/mGw8sVObh7jzoHRaKHumEsGCNRQKMZMmqrCyLuYTCY6Qp/jpl0hJhbF/3+s0hRMK/
qX0Z+KSfxdtUzeGv7LRUqxxwAlO+O9T4ue9joaTGZHPtvgraAQHZMck4aUH1d5xW3voGjckAN94r
qGiFCz5In4KSw3Xe9/Z5vvI+82Hn6uelMZpw9JgGYWtEcqrej9G82K8SRNxyBhilTuMsLYZY6lk4
U7XmBeMT5IecUHSLsOxkgnMgYWe6EmjawoZ8SIOhT8YQ65X545crafL9yiH8DuKpb3rGDOLBD3/7
1kgFfv0GpQXC4eXgtLCLararjYNX6bkTMYbzl6YJscJXOOCY7NxVSbewdEi3ce+bqU4kSqLGK4qK
kYsxPtXhtLjOvfgReBdHE2+5O0kpIGUqWgIi7As4TvCr8D/1teAo9Zf0ww10rBT7cIbuDxMGDzMM
xt4ln97Ju56YFDsIWAOeukFGELUsspXVERW+6J/F0sVeLiqP8QGM3wutY9azaFcPv8OP6n8xmIFa
NUrbU/NQgAv3amz7iGeaq7ZDVb6zIke3WnmlyHWmeVNi71QMbpKNc/Q5JXodC/539YOtPZ45odwQ
fItcYG5SlrqXsTkGNH7/mVsB9+DlWsZIB1ID1j5n9Xja7E/W5WLgZiV+IfNiYYlKIuRtAWeZzVA9
ITONxNeaM8yxLZQlvJrbUuJGuFbK+8i6Z5VqnfidWgo3/q8I0n00w76N+X02whde/xwUFFW2Ojdt
dKsOz4YJT4aVvKP4uuh+0nCqyUvhKU8iUmPh9TmJm5BDSko/+vJ0XTbyDOmZ1+V92ILbDRnbrveg
V7KC+K81iRuE3T3vu1ZZSbF/kXr82YubzW7qcuZpNtBeQRyRqHADnHN5o8tlAEF8xSIv81Rq35Uk
klL++rVT6IksWQVdtMlipLW2ZkaARz3cksCZZTzbCf5T+/feLFE2M+KzeD+ElgVlht4dsK5muEiD
8zIGfUN+MdbZrajf7XLWVhCDM31FhaqmvNb/GayyCKqnWO0OZ7z9Ec8GQXIspwvRLt4Ug5NHveGQ
JVXVVUr/nGEyPwH/w8kkEnrSXkvO775muZmwL7I7vuLScf7jX52B0hpCKBjDZvjFsBMXsy+7veVI
t7J1fh9VUh8fWcnAw5BBu04ohkrOrFBOmXkpA/exkpznkjkBNGdxI4H7qJRZsgCIMMC0g9EThskp
nwVb0DQ0i/mMZC40sU7wjgdtSQ2YaieqgT0nBSSYrwpcoDgvlxN2yLfOdXc/S7RnaTyTFAL15TDh
jZn8CQizaFWVQrUVYE7HP4BiPpdQd0j7vAqt/S6LBAmQH9x8CO8vTxUQOXLhcTctP7IyfJP0SXAp
5lV2RlV78r/GMbYgB+aoXfQ+baynuDmU9nHgkssFlRaDjWDJAO8pWqLAVRyP6n0k/T/vE4JYyHva
aXe1k5PDUulLfaPQViAVNnN/ojQs3XTjhVdl9wIDvUVfw/3HugYGpBpwXprCwfBMIM5sT3Eohpzn
v/Ij9GkyvCbwfrS+b4pYFwFvS/sn+U0CDrScAHk3RSdEQgJnCyOboRdZ4cOY+PRD9T64FTvOFwty
qewAn9/BSB5VolnTabxPxa9p2JXj8sJ0T8cXfIYWipo8nbIAFT1sSWdsQiq9pzdzDxv0VioAiXpx
UigWxfT6bnH/ubd6ZnFmLX11XsEhRSN0DmXdZCvZ262d3XM9V662Qk0XXXfLJUo5HzNXcOsNEJ42
8O5jaCaZb71jUvoxv4fh6rZrgDN+dB1OAfw3zejCPUTmT5/QLtHd9POZmJbO5P5BoZbzyg7plYMR
qfI3Sm+SkBZNqnjffyarFqowsNcS4OlKuO3OVQCSsGDFJ4ePAhP7n1xYhNTY2ztweD/aeFJWmQGW
+fmMySb7wqZELKiw7m074yC17qNYyulOwAAAmxXJybP5sBv3hraWb69dkzdc5KmlqCoRe1eIrmBv
EJA820EOhpSTm4XUtLpOrPlWAux9mNotGaq5rCnpUF4TuSpIJtyRy88iitl2VYRGKap9jMFiTzQ7
vPJlHH7+4cJWHA448RERfWuHbHQaP9mvgyIgMaP3SCK4Q9QYahcPr/Bo6DeU+XMrt/GGRutXlRuf
MHiqtPEFf5kA5kL//L9p5xKL7QBZ40+XdMyFkhZxLgBjfQdDXzL37siMTc54BSeKLzh0UY5wtmit
jppWpply0tLm7vRiQgakK2P6reW6WJKXQ0Ezrq7yw85+iHv6xWYv+p8V1TprP3Gd0QdmcyVAP1tC
DMdb5YFLjJsXVj6EbcCVJ/BrjEHg6BU3drBcl5CD1APAKoxtSKcNh5BwIF57Bw2Phvu2A8ZHbvoz
qfmMZdOTMLJ3WpfGt7XfmY1plz8H6RkZFR4+yDE7IjacJQvy5S311cNgDi7u170N3x4Ik4Ibeqoa
AgoysE2dDguY57Gj5pFJERrIKvcJNtTZhOPQ5RHhjJPps6Akyf/Bdi2lz1AVZzB8hT9c6BZit/bG
GKSXKqw8DQOlTnyX+NeSuB9BOhp97FhNZu42mBzBXmLWNs0DceaHAKobsQH1i21MESi2gArEm18o
kged5i52IbJsk55YhWulw1xLIqWlgrpecYKD8l6jm721Eu5aV+Aazh4L8jWbtyrsfUKtXl6mLrgv
9HilGe/wp0wgNUDs1YxhoVMDj7P8thClAGqC7puFnmXERklFJq6sy002FNQ/ptIubwFEfxFHJXPg
VsDUbI09h357E8rNHFQTn27Gf+yn8JLEweUWG0O8Zs6cF1eWNnEsUs2CtOvbCXtgEQK3oiO9BdXH
165/PAnsYrGAcozmPLFLmpEOZ2WmghYuj6w37mtLEDOFiVWplsMxhb2wLgJiRumzCY/v2lZecGLq
3939kSXyqqGgF1pxRfWfc/mVrEsqLH8KcByZLYjgTucZVLbfo9QjuwmYup5JEn4Rdxy3XVEJ+EiX
pmTxVoDskcI8XWRzdxdXcbDyjvGkg4GtMB5afOiTuRKO9KRtfMy6ONuXM+DK+H13E62Quy6ldxc8
cP+eanyU3ulOZHrp5tJCeynvbiMADmbemqb0rtvMuac8mXJAXoRoT/vH1IUIK3s1PaPzOAUkZzrt
rZkfYo11dKglkwfwi5PcktTLjvNEGZIs5dmUoycWZFZ8MTUz5ozZfeHE8tzvvwywqVTbTyClgkIM
6IAsxWhDgeMF7fmh2bLnG2oJ5nVYDitTdjLtd28llS+KReWE8zYLA43sIAsa67mf/IbDxKxcAZmk
fwYwpRhCtyYOs8iM2xNH1FBDn+P12hIgHZEJBLLczA9brua4tE3jiUcNGmpf6JIDkrwdso3SlB6e
IxLG1QyQzF9Ax93IRaAsFbdn/chdObcjxOXc0yy8Qk4PZ192hsmFWBZF9xNjro9cCgQGEI4LPn32
K2KBkPy1oVPMSLMOs+UFOYElsdj/p3RlY4bdRlFf6bkEWB0AYpIOuaa6arWbxDiUmjvApP2WJ70l
f6KXturfCPRKQMKvw/sIL+9i7vSobQ4tzxGruQlOoR/kWgJ1rLuG0dQWBg0ea5ghSqCsRfX1xUtc
gFKqj7fvMEIHJjbmiAaanpAwON02zljvSTggLCRxxInN/U6HSXUnA1c74o1K5T7TI60HgoIGIMai
+Pa6+Hvt/Jr33a0sVBlKpvdcCLBmsBP40YdPGWg+ZzquDI+nPVZ3gxdBMa/dVtOk03z5eihYyKNh
mjGLYZSzJHTNL3Hi5XrLtfmWG3ak31bY0Ec1B4PFrPDbdf18SyMycmGcgEfqcXLOtKPd9A+bVS1C
tEu9pUMufRFZTzcPH8FbNwN+E8F/WPKjPweL4TjSYqSAAqGxGUcvu2gML/k2WDwyOnRHWODMJ+Ct
ZrmfAnCbaKjOMCNTjupTQD09UEvCjHnSIBu5uWEAhIfuRZSnkjh9GkGFIDeYCrL7WQHwGlcFFPDm
9vCbIPYDK0FKAx+QdQ+tffyTLtgz95yTmuNukFjOd0n8qfU7f9jo3aoV0k2+BFfEqE9hc/FXi20+
kFuNaqGmmnfzwZAVt75IjL2MR0YLO2oE35LYwxEw0vzJ3UtZhF8XPoriPFmxy24AekiMgvReFbNr
V71e5P5SOT4OBio80lBNz0ohIf85nlDWmOhWcb92yQLgQ4NTHcB5Um7C1EBXUG/KeQkJ7LHzKlzO
ujuydQU/q0jJgYJif6F1746SsergRIifOTMRqFctPSNgRg2u+ew+Rl4pW0ZOHqe0P891SMeDUQEX
cIXcq5BaZeioKN8RtJUPfAe8SDH4oorEEv4IM4LWBiDFEY22Ib7OvxPLP4zlBxFZv/JWl33E9Op2
cHQG8ABl6CLYQgVIYXp4kWvpsehfRcQy8AyXvALF9hVpwbQ10hoakQW+3paWGzfTngPqDgBfslN+
6IM2UqNMNnatvnHPVyIQYY+B7B/IFHAuF/2kgIb+YBunPew5lEr2ZRBfgz4XFfLyvJEGlZB+hvcn
LGFerXR5QgMlSAsMuqAGfg5tB4Ya3zeE2Sso7JnOGomM0eBpBeSE0GhQRl0foV1rgnGZXqAiaMjz
WbgyQ3025gRpl2hP8YNc11nMI6UK5VE6qulx2mWQJyWZtXYESac+qxsMCO2iKFUjVyZR6Cln2f43
snn6T0z+ecJ1P5J92vWItRuBMh2zAmAonFQo6eiWTyguWUs98WewXlOovLCdXULHKbwvZjq4lVjx
CJ+ImxCPv9t4wMCr6LHYduam5OwxFeKf06/VSyVZToNYLUN6DHKrBsE1I9sKWUI9B7WTOSWUDpgD
1YA21Mpo1bUtz0XSXab55aMsTUyl1OlCy92HOzSbCeVeBo5Id03VdKOimXfOnrAsToRd2rkleha4
UchYrxz+9wcUQXo3fZn8xCwBSvE6mShgNN9rYLx53v5yjcU4069AII70HEK6SOvNCnim1NQ4UxXP
N2lIZt/zDF6dstL7YQGAgwiYMQdiIomCwZEKrh0Fpic+mUjjWMhnMr1REUkvZLvjDph8bo8WRHwh
43ocbI/2o4nvEvn8p5RJifElHJpYDKBeAk0/tM1nFuFKpTw5Crm2yL45nHcqGL+AgFeSEhNh47O9
AaIFFeVxpjPiuzbKz8Y5MdlEIop+QwAAR/RasxGhSQYcFtIjHR2Wizf87UNBj/5/YePgsJ8l14ZL
3xfdhHynLZgTZov7No1RTVxbFGo7mwpf5R1hyjDte/QgwP9qus5Awt7XpoQyz+h1EwVkbqxVySO0
HscbkzokcFhX8XVgWnX3xJo3
`pragma protect end_protected
