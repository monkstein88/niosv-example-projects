// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
TvFlfTOSkk4dTXM1o+DTqniW7xARvJevBKTkJN6HdzvnIawbB8D/+dMBC1vfPHt1iQSqu2vRmpV8
cdH9p5mnadCbwQm9eb5hB2nOJo2phGNLI3n17UTgNJq1yibUGP7b2hbMFeoGlkg4/GZBIXFBvWXw
kn673JWmzuCfZK/Ycu/BtgTWY4X3Xwzzsx0p4wZJZBGEJOr2cftGTBV0ebDcsCTcINEZj6johHdB
63ks+mKqk+N73MptVQ3lvXAYRCf0VTNZ5MEJXw89wJzBUmJ0RWvv3K91OUNzQJ7++FNuKXfIMwVJ
6p6ae4lcPFe5LBUE9sQD+aNqyPzszAKdeR7OKg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5328)
iSqPORXP9stLDq0MYCjmZETTHm/kje5ieLGNBApGWCWb5aVWMyaUtT5sTbf7qqwgbY+yid9iYBav
sNcroI3LOeDd123YVTPoWlzRUz5z11BEX3Pz70PQbu4nY82Jc4+5xTCu+4S+dyPtvLgybSDOlU7J
6Y0P0AVQzsrg64gaIUp5f6WuEWc6jgbCz3FYPeXBtl9CK8Yk4GmpM5TsAMAYstAY+QoWWBiOj5xX
mrweS+ieg0sy3QqyG1M2yrJLOHUliPNKmUjL8msPHbhPL4gPeuehQxr/FgE3V/U2NHuiHI0DCVVA
HUAB7WhX/NqQhOY6of04YVAb7cx8d7qapBr382WHfoRKivMtPHRQCMAS85F0HaTR6YiAEXJjktmr
AOTKN3hzblt6uF+Onda6qMggoBolKYhTg08PzQ3RLoyAmAcsuw6UOV71ju/TKyEHikc3Za4TE4oy
m6mDq55tng1ohKI97J+I8hwVbVLzGI+ZBQvxoXhaaR9+bB6+tBDLrMGYnyfE6lY0XQGqYvAlZIDz
E0vfyzgafOAFXPzWCMcT6L4uORyJ/I7Qi/UB4hBrVah9+YdCYgePkuQO6hBAKylco3rceU9bTgPz
9Ynk1/FnI18jyfXZEsrFJNnxysPwXKeeNtU0GB7DK5wZu8QoySyIJ10htzEhSfzn0A45pxcq19FB
dIIXe3Naa8hDkVcRjh4Nx3R0UIhEnZEPVEhT1Y58R7KetuEW3Hh95mZN+pYmZXBYl0jsgeXPWhD2
ZXZ5gDqsaTmmZPkynEs6CaR0/5Nd5PnbV7Lp1nXq8A6cXbgi38fBhONUT2ZCE2t5O8dP6Sb7GdKc
QVLmQzg1ocpOULM3ga5xQ+axlufljX+PZefpO4bbvO4BvQNbG84BMiBZ8tAItUC9cYXMe/zbarPJ
oEzIC2oVqpwvLm3U/H4Zhp6Ad3WahxNZ+GC6w4/w8oohVEOHFoMDXE1+n8hN+6Gw+fV2ikzjB9mp
2mbHJf3OCyhsonLLQvgeonDgk2jNLbXKF6u3RQwKIhGoLGANxGhT6gsKVlCEzC6gvzZZlRdmEbhf
bVBD1hDiUwg7Isoo4tkFaGQG4cKbODO4mI+efbEB+ps72NOCwCwab1ej3GqPQlMtkxzMQwDaXcgv
zCw+BhX35msPxAJPOSO0gicJLUCWF+nmWxGg6r1SQXGpRRzSGZa7CxVVO+LcgP9/O/rsaNrmVUtk
aKwB+ZE6Ltekd6juGWCwV7ZNxuV7fgCW0GcSfCA03pn7NQZWcJQByJFWRbCEbiIKxb4f6b8Y/cDJ
uIlXY1aYXy2Sl6Fr0tuI3mSZi9YGjvVG9BoD8VYR/zDLuEBUz2dJ2S3zCsVVkxOX+p7pFoIAFPai
cqf3cCe9HC9ROVo2ajUYlB29SAEb8vhbvSCp0bErLVkt+24A0Wj4topJAVgyehIGrVShvw0ie8R5
32FjDIuvUjJoqHRmcwJc7lSqN4HS50I6tYpyvq80CIpMq6nT8uwJ9HEDJHj5CTtu6eotEOid3sXS
W39jypiL2cH0FCfJqcNGg3E4NmDv9vOJVSjKfpfmWQGKIzI6yv0RCFx1KWpYOiY9Da2ERtZwIn2K
nWwMg2jHaw9nWWeb2rzhU4Fj3wiOm4As18Md6iVEP7bS/kVlmwp69q2rIsY76YvDv7R1mUG2m9Pw
gC4NgTzQmVgGMxoqf2s0cW5P/7NDVEVC2jKK6hrbfmjoS6FoErmlEZqNXXItLsvXou4fSJFEsp+v
1bgVSynOTKZ0xkqc+wYVuZ//x77mB5meduUbCQmzrQJm50Pe1DTkgtl4U/MKuLdaz0KBZKEhQ0n0
22BXTlbbT7YQKCmNO7md7trrXs/2eB5qCNOdabH33ce5URS11PpzZWapH7M3xBeoWnWxvtfnrT+M
dXIrg0LyBOAcO/Zw89btAtes8VtyYWr21ckOnPUt1pFCMOoSa0NeN2ffcvcBNSQ+MRHwGN2csR1D
cDZimXDJS/PgN2fXHK5+d+xfXLtdC77jrjvLbJA1SqG+/QDZcZwzFnY8IVEBCJ3qqq/jcuYRV8ey
U+iWE8H3gHCdVIS8K7sJhqSzHMR1jeID6RTXZPKmGpt/OW9i3R2sJ0yTfHImp5OjYMDAGdPQ86NM
HZJJoigcMP3T2uMgKFSG32vIiRKvxzgTuQB//IxVVdjFc41UjCKFsY73ZePq1GDV/NbYJrX7a23B
YYirlcslgEJMjNFR5Aw9t5Zrv5jdGBijWhEGgMKVMKCrJ8fN2pa0+ruGvpV667nd4ALlsp6KyZEy
q4rjo+evnQt/XB5K4CnE2SV4PJrppISMv+pQ1LRjjERo4nuEyk2syyfk/KdWi5AQHz9DZBtl/Whw
hW8PlQK/pZ9EeIKfTf5UTInRc+B3M1IjJoITr8jsamBiPM7189rN6Kg49ghY9vrdoWaOO95JsC3R
8Ln90mAo4hVLBZxarOu0pEQPOQT0BQTkugWIkMlShyVevc7kcUPiyMNsmRxicRbIXZLhd2pvIqZJ
kjueWXd2586dhbFZw+kvEmPHRtgY91IXR2rGxrIjf7KFLN9bhz2SdWJzQ3K3Dp1pAb/pmip1ihMq
95nL78SxKiMugtV2OzAO2bMwjG/jqA5kz7JYEnPS2zy1mdD0dIAoKbQHTmL2QcJz9Fw56F6lD2hU
f+p0fZIKpTnIRmBhTZSxUO/0QVzhKUXvKy2NYMiKzSPhKD4vn4Cr+j28NvAp27m4GZxZHE8UBaht
md/yD2L3Tv331LOjQ40Ir/Zc8kD9KTEbkEZEOx6uUJfmMz2/r0WqYEmBBfam2cNJ9W/RjUrLk+sB
6awaELODhYGTUVaqjP+1vChHQ9hgQ9fLhpGc+cAFMZZ+seADNixcJ0u2SQrfh961blpTX2MhkSkO
+8nHzUTrVt8SK/4Rq4OewPV9fAqWA5iCDo67E+zuSFbXmNKr58v77GdYYOPXhsf4M+QNmJ/s5nyd
KFDzpyusEKhS/EOnP3WE7mCP2Lt/MA6dfqq5SxTdkX3yUZ0kxdKRNjxugOfp9bRgGCazVbgoXVre
+dT8GWeY4RGBTT7oINURg3bd4uWfz0uq+tp/rcKo3jtCbYvmjkXrW2IWTqdsCVvrpoHqOAYpZ32k
BHk/ey7aTIUcockAbcV9pnQpGj1dfVeqkFiPu+LdUkXFE7VoeVb3aK2ouZTbdgE6il3TSHjrt1t7
jymaXthGYYh7dELbfCSy6UB2/9izOd4kvqDjINq0EXus4wOXDwb4DpF1+eWOF/Qy0xAJTtFETbHm
dO0e/pMraTf2gV8HFZT1dAZGk2JXKb/1EzYUx39X4U1DFYvRC97u5JcZvOePHjU+XZzxg/1y5Eb7
xeGQwF3QwN4a4Q/I+zKHcOz29GEk/vvbw7n415Nawr3Bqe6SFixkK6//9Iri29NgyQgP4L/rGrAz
KlsF4ynumJOTdsu2WcZUTcExJkxkEq38wks/TaF8q7ERw0ZMHIS4qi5YA/8FllPHPxKixFrNLfQ2
+T4b426Vt1LVwhKOhbl3SqTYtcUJNuuMC8otOB/uOp6GCDlfv6f8wOVZu0rW9mwx03BebTpzyflc
XI/WuLbCONVqbSkj9r4p+F9ChATR/owC04Q/lMMXq2wQgY2aJiCeGvzNEDkuNw4utP5ej7nSZ9/l
eVvNbATmk7w2VjCfgcRmaDCXpcYt8lZmnh0ooY7fJzxXVPh4majmI0+jEvrwNjJvxOAWSt+M1+4v
/fMP6XarLFAWBGIQDCJX5/3SylWEycz3foIcJmkYQBkN9DjxIgravD/M/JgYznkzWLqtYxxokfo3
sPwFzzuncQ0gt6gseimZQQO7JC1Wxuvxn4bPDOIGcFZFSxmhXpPMvh9Dq974cU32jFR0npCErU4x
IrebySiYiNUAFgJuU/7TuaXNTOq0yIOsaB1RNEIU3WxNUl5+Lkbao3oQuJgLSrnvf/osomlu+PYT
2cZlATXrqtfm+y8wJqifzBmeK+/K3ua3P2IyGF6Pyc3NuufwuVxQUnkLX/GecVVpBieOzMZwFUR8
3mKhgk7Rj0hYDBXyNespPVx3Faj/3MmXFaJ6A00SdLY7yxuaG6Is7STAyRDfPD4JTMzmpXEfAehk
HpazT63UBqfriRKHWmM7iLZezL+tJLLLl06jy682Kb1nbcZBGvTdAJWWNgJWP/lGi3UgxrWPskk7
RUWed6fG4s2N1bLonEbaoPbB7IzcY/fcpgRGLKCu9vEnNJxJS9Sjje+RaxACRscSlfSLL52IBMuU
4jvaXt6j+88fWyQOB9YmlK+WGJ6983AEjZs/aFFYCiNTvO8SyRcDSvxjoA0ZMs2qcwKsjJLwJR86
tYzwSP3MXLnXHtuvWmTIU3ZWvlIDR20RBKWT2pyMtDpXqwjOmFeRQN5guTdP5NEB37dx2pX+24Ri
aWXrYE0s6zSsYsQ8uJWb+fVAjx4Fu5Ko0HChLPwv3M57LY5CbzQWJJkm84CzCaVHXPq6BchZz62N
zwLjDNDthrLUYyzalg6k7ASUgC/FNcjDj3IeZpQntmXtNKJkDD/FC+paE5ehMHnDgh4DDyc4y+1R
lfpljbDi5BD51uYxVEFFGvEjVx37wx3sWoNbfk0Y0abLj2+0CjiE6qMr5f+BKBWeTTaBac1shg5Q
RybV0p2MOobUzLl1SLhZK6yyQoyo/IUIzvnLdywilQ0w4ZAwDDPChsAwfG3qZTi4Kahxcr0L4u4m
OP3rtNA3/aNQpGcnQPKE+bF7Sb310ohxmSoCTWiJ6TyZDk5+a43gcyztLRcod9rxbMMhqbDIczS9
3ZK6s6uTG2SGqD2esyjGpROWb1enjwo3Zb875KTw5X9o/jaqwPrPkm6yOQWw+8EQ8Xxa1l1+7R6t
qsVJbTNkDqbHbylAr/5CcmhDrNIeduhcnYJRrT7rTRnDAupEraDE5u6orOdwCh3R6ky9p+OAMGT/
uXokNXsteeOaR/8XkUSNjgmIOQUEbUDCpb0t/E5dJqZd5cVTLbYCORzyNL8dXi9geRGydHJbPFSY
oN+59z+extFiS8Xe3+RdHk4J5dUlGj6dlSQ/UY4A/bTUPjBB+zzbsEfiDInSLZUz7v4xb3iAKw7Y
3GzBwz4p8rumTSfsog3RXfM6cXHs+Gg6hKqeI/hKBvszTZoigHxymdwi+uDIIFCKHfckjUpc5IjG
nhs9G62bYX0uT82dRqseMuhiLI2xsnv0vdgwGNhFZffInU9qB1fecuS9cxFFNcCoxs4Ra4nP6Ypr
PGs1XSZfY09DUyc0wlR5qryVHDe1xA90NnYa9Jtns6hXs5ppA5bu7FslqB3H4tZlT0BhLeEn8yuH
BKJGnimr7owBIZZQ76cK14nCBKKiBVwZTDlJSIDSDgDNQvhvU2SGV430OaUux76HmcMdyTxu1/vO
ms40h74Foepm8ieHyO/WuAcRDf9TEo4fhD9muMBV+tn3pvjp6rgMOwb5fzkE3VbXHgiAnC9GnUYu
GVtrJgySH1u+NGv7AZ0TszDmxqxO116iHjq4ha+H+NkExtdDdoBrdGtrfKLMSaQ3pHsftQW3Osyp
7pbIRdbtE6z4r5z3w4TvBgxnUDJqFXqoK0m+OFjP3KBCKEr4TWLXVPVeA6InuK2B4uGLFqDa5sxx
bh2GDYD9TJtdFOOxNaeNSKCTGx6KXPbS3PAIKoFDFddFyzty0oyinZolnOp05jTnk8YSUTBu8M6Y
2MGJPA2CKkieGbzEHDjE3E1TNYRRayZdI+CrIvz/8/Jji9zCaWWfi1euEqrP3vdheeHcsrmj8mRC
Qlde5Y2/JFh6+0tN6M8N7t2AKgxkJv6JzhPSp2DYVYYveV3NctDCTndU/FhNUZfPIq5pibZR5UTZ
OsiM23uLxXDXFlhmPmZRo2mHrcG5h4UK+HWDt0n91GEt59mba5/B2AY8iFBHVFLjDeIkWj1uR2Y2
IdAzvR5X+qS1v1e09l2POqJZWEaovpK+ejlf43NBOyz9lzqCzNkY50boIjwGNei73KriUdm5+R4A
CA3beNDMQuCyARJYx12iydn5tRrraIw/t+ZZEjUiePq/tDy/tnpVu4/56XnehU/sae/R8ImIQHak
4XqeO9QsCVK+HFUdrfm8zOl0FLPR7xb1FL2AoiB9waqzWOifEHiHbv+eLLh5aMpvO2+3sTepUazT
E1693s//F5CVFPe+T89Is/h0ARgo0ZUXk+mOhIRugQWIwgcvhueTD0Dj9+T0LE99T+2njdcKFi2O
L9/r5IA7Fzln7L8XzLWGZWMbrNdi/8+xb6UjUv/WqbSfgbOXno6EFUmsy73wlD46ih/9jv1B+hlm
kEulC2tnCUC3mHR1ptIyegKcaWEjPwSKfqB2lw/rNGjexJL6mQijQzD6HLQMh0+IjGB2NppQRVxc
SIS1rmJukhBbMpPNOU4qQGQs7Ef87rfsPk1XmL2jj7t1r7UfKfTyPERW8TCqFroKxwG6UHWsEdtN
L2SUfTM/IZDSu6i4tKPLY+6SpH/v4R3MhHAGJUtyZCGj3j8hOGf3xgf9oaM8NcCy6zcqw6ZFdsVd
/hVrwIGHruxQGbVpi9dlQFkNGU7WR+qjhgP56QWg7SNfVHyXefxPEawqMmGyhsJvYQOjJ54YrCa2
1ia9TPzCgMxnTdACPMJ2sfxIG7aRLDQ11bmLbMVMlJVcGYQN8QT1tRyMWVt5jg3HIOQ1IDe9XShA
kgt+0RpJqoTGoHJimKEZzZZf2eiUaSQdE+7tlU4wnjLvBHMxwjIP2omVOIWYUxRgNG9zTI9uSt4D
QdWA1Y5CehIv2zxgvjS+SuvDl3aT+TNYxImoNu8I7iPfav+Q6LJyMTHyaxbBiI9zQuhBlMBIjAxC
3d4qaaLx/s63X8bkiUr1rt+OfRldGLQjTpzLl/WCAzPSE/C5Iq9r7I50b7AcUn6C5ddU5td169ia
RC0JuCU8FnprvgnUakvNgftVYV37BP1KNREjxkd2MZJmdExPxzD2KJ+QjvpjmWlIkV7pOHSrGwKM
97rouDi+61VqJ6xFQwPj5B6u0ChmUpBaISBMeCTHpnTp2/C5wW+qdqOqFKM3dcRkLmIZpaFgkxgm
q/4H50/Jo1SA9Mf9cSeyP5DyUdqOCwxioSeG
`pragma protect end_protected
