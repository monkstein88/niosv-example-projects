// NIOSV_SOC.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module NIOSV_SOC (
		input  wire       gpi0_butn_external_connection_export,    //       gpi0_butn_external_connection.export
		input  wire [3:0] gpi1_dipsw_external_connection_export,   //      gpi1_dipsw_external_connection.export
		output wire [7:0] gpo2_ledg_external_connection_export,    //       gpo2_ledg_external_connection.export
		input  wire       in_clock_bridge_in_clk_clk,              //              in_clock_bridge_in_clk.clk
		input  wire       in_reset_bridge_in_reset_reset_n,        //            in_reset_bridge_in_reset.reset_n
		input  wire       uart_serial_com_external_connection_rxd, // uart_serial_com_external_connection.rxd
		output wire       uart_serial_com_external_connection_txd  //                                    .txd
	);

	wire  [31:0] niosv_m_cpu_data_manager_awaddr;                               // NIOSV_M_CPU:data_manager_awaddr -> mm_interconnect_0:NIOSV_M_CPU_data_manager_awaddr
	wire   [1:0] niosv_m_cpu_data_manager_bresp;                                // mm_interconnect_0:NIOSV_M_CPU_data_manager_bresp -> NIOSV_M_CPU:data_manager_bresp
	wire         niosv_m_cpu_data_manager_arready;                              // mm_interconnect_0:NIOSV_M_CPU_data_manager_arready -> NIOSV_M_CPU:data_manager_arready
	wire  [31:0] niosv_m_cpu_data_manager_rdata;                                // mm_interconnect_0:NIOSV_M_CPU_data_manager_rdata -> NIOSV_M_CPU:data_manager_rdata
	wire   [3:0] niosv_m_cpu_data_manager_wstrb;                                // NIOSV_M_CPU:data_manager_wstrb -> mm_interconnect_0:NIOSV_M_CPU_data_manager_wstrb
	wire         niosv_m_cpu_data_manager_wready;                               // mm_interconnect_0:NIOSV_M_CPU_data_manager_wready -> NIOSV_M_CPU:data_manager_wready
	wire         niosv_m_cpu_data_manager_awready;                              // mm_interconnect_0:NIOSV_M_CPU_data_manager_awready -> NIOSV_M_CPU:data_manager_awready
	wire         niosv_m_cpu_data_manager_rready;                               // NIOSV_M_CPU:data_manager_rready -> mm_interconnect_0:NIOSV_M_CPU_data_manager_rready
	wire         niosv_m_cpu_data_manager_bready;                               // NIOSV_M_CPU:data_manager_bready -> mm_interconnect_0:NIOSV_M_CPU_data_manager_bready
	wire         niosv_m_cpu_data_manager_wvalid;                               // NIOSV_M_CPU:data_manager_wvalid -> mm_interconnect_0:NIOSV_M_CPU_data_manager_wvalid
	wire  [31:0] niosv_m_cpu_data_manager_araddr;                               // NIOSV_M_CPU:data_manager_araddr -> mm_interconnect_0:NIOSV_M_CPU_data_manager_araddr
	wire   [2:0] niosv_m_cpu_data_manager_arprot;                               // NIOSV_M_CPU:data_manager_arprot -> mm_interconnect_0:NIOSV_M_CPU_data_manager_arprot
	wire   [1:0] niosv_m_cpu_data_manager_rresp;                                // mm_interconnect_0:NIOSV_M_CPU_data_manager_rresp -> NIOSV_M_CPU:data_manager_rresp
	wire   [2:0] niosv_m_cpu_data_manager_awprot;                               // NIOSV_M_CPU:data_manager_awprot -> mm_interconnect_0:NIOSV_M_CPU_data_manager_awprot
	wire  [31:0] niosv_m_cpu_data_manager_wdata;                                // NIOSV_M_CPU:data_manager_wdata -> mm_interconnect_0:NIOSV_M_CPU_data_manager_wdata
	wire         niosv_m_cpu_data_manager_arvalid;                              // NIOSV_M_CPU:data_manager_arvalid -> mm_interconnect_0:NIOSV_M_CPU_data_manager_arvalid
	wire         niosv_m_cpu_data_manager_bvalid;                               // mm_interconnect_0:NIOSV_M_CPU_data_manager_bvalid -> NIOSV_M_CPU:data_manager_bvalid
	wire         niosv_m_cpu_data_manager_awvalid;                              // NIOSV_M_CPU:data_manager_awvalid -> mm_interconnect_0:NIOSV_M_CPU_data_manager_awvalid
	wire         niosv_m_cpu_data_manager_rvalid;                               // mm_interconnect_0:NIOSV_M_CPU_data_manager_rvalid -> NIOSV_M_CPU:data_manager_rvalid
	wire  [31:0] niosv_m_cpu_instruction_manager_awaddr;                        // NIOSV_M_CPU:instruction_manager_awaddr -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_awaddr
	wire   [1:0] niosv_m_cpu_instruction_manager_bresp;                         // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_bresp -> NIOSV_M_CPU:instruction_manager_bresp
	wire         niosv_m_cpu_instruction_manager_arready;                       // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_arready -> NIOSV_M_CPU:instruction_manager_arready
	wire  [31:0] niosv_m_cpu_instruction_manager_rdata;                         // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_rdata -> NIOSV_M_CPU:instruction_manager_rdata
	wire   [3:0] niosv_m_cpu_instruction_manager_wstrb;                         // NIOSV_M_CPU:instruction_manager_wstrb -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_wstrb
	wire         niosv_m_cpu_instruction_manager_wready;                        // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_wready -> NIOSV_M_CPU:instruction_manager_wready
	wire         niosv_m_cpu_instruction_manager_awready;                       // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_awready -> NIOSV_M_CPU:instruction_manager_awready
	wire         niosv_m_cpu_instruction_manager_rready;                        // NIOSV_M_CPU:instruction_manager_rready -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_rready
	wire         niosv_m_cpu_instruction_manager_bready;                        // NIOSV_M_CPU:instruction_manager_bready -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_bready
	wire         niosv_m_cpu_instruction_manager_wvalid;                        // NIOSV_M_CPU:instruction_manager_wvalid -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_wvalid
	wire  [31:0] niosv_m_cpu_instruction_manager_araddr;                        // NIOSV_M_CPU:instruction_manager_araddr -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_araddr
	wire   [2:0] niosv_m_cpu_instruction_manager_arprot;                        // NIOSV_M_CPU:instruction_manager_arprot -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_arprot
	wire   [1:0] niosv_m_cpu_instruction_manager_rresp;                         // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_rresp -> NIOSV_M_CPU:instruction_manager_rresp
	wire   [2:0] niosv_m_cpu_instruction_manager_awprot;                        // NIOSV_M_CPU:instruction_manager_awprot -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_awprot
	wire  [31:0] niosv_m_cpu_instruction_manager_wdata;                         // NIOSV_M_CPU:instruction_manager_wdata -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_wdata
	wire         niosv_m_cpu_instruction_manager_arvalid;                       // NIOSV_M_CPU:instruction_manager_arvalid -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_arvalid
	wire         niosv_m_cpu_instruction_manager_bvalid;                        // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_bvalid -> NIOSV_M_CPU:instruction_manager_bvalid
	wire         niosv_m_cpu_instruction_manager_awvalid;                       // NIOSV_M_CPU:instruction_manager_awvalid -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_awvalid
	wire         niosv_m_cpu_instruction_manager_rvalid;                        // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_rvalid -> NIOSV_M_CPU:instruction_manager_rvalid
	wire         mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_chipselect -> JTAG_UART_DBG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_readdata;    // JTAG_UART_DBG:av_readdata -> mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_waitrequest; // JTAG_UART_DBG:av_waitrequest -> mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_address -> JTAG_UART_DBG:av_address
	wire         mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_read -> JTAG_UART_DBG:av_read_n
	wire         mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_write -> JTAG_UART_DBG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_writedata -> JTAG_UART_DBG:av_writedata
	wire  [31:0] mm_interconnect_0_soc_sysid_control_slave_readdata;            // SOC_SYSID:readdata -> mm_interconnect_0:SOC_SYSID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_soc_sysid_control_slave_address;             // mm_interconnect_0:SOC_SYSID_control_slave_address -> SOC_SYSID:address
	wire  [31:0] mm_interconnect_0_niosv_m_cpu_dm_agent_readdata;               // NIOSV_M_CPU:dm_agent_readdata -> mm_interconnect_0:NIOSV_M_CPU_dm_agent_readdata
	wire         mm_interconnect_0_niosv_m_cpu_dm_agent_waitrequest;            // NIOSV_M_CPU:dm_agent_waitrequest -> mm_interconnect_0:NIOSV_M_CPU_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_niosv_m_cpu_dm_agent_address;                // mm_interconnect_0:NIOSV_M_CPU_dm_agent_address -> NIOSV_M_CPU:dm_agent_address
	wire         mm_interconnect_0_niosv_m_cpu_dm_agent_read;                   // mm_interconnect_0:NIOSV_M_CPU_dm_agent_read -> NIOSV_M_CPU:dm_agent_read
	wire         mm_interconnect_0_niosv_m_cpu_dm_agent_readdatavalid;          // NIOSV_M_CPU:dm_agent_readdatavalid -> mm_interconnect_0:NIOSV_M_CPU_dm_agent_readdatavalid
	wire         mm_interconnect_0_niosv_m_cpu_dm_agent_write;                  // mm_interconnect_0:NIOSV_M_CPU_dm_agent_write -> NIOSV_M_CPU:dm_agent_write
	wire  [31:0] mm_interconnect_0_niosv_m_cpu_dm_agent_writedata;              // mm_interconnect_0:NIOSV_M_CPU_dm_agent_writedata -> NIOSV_M_CPU:dm_agent_writedata
	wire         mm_interconnect_0_uart_serial_com_s1_chipselect;               // mm_interconnect_0:UART_SERIAL_COM_s1_chipselect -> UART_SERIAL_COM:chipselect
	wire  [15:0] mm_interconnect_0_uart_serial_com_s1_readdata;                 // UART_SERIAL_COM:readdata -> mm_interconnect_0:UART_SERIAL_COM_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_serial_com_s1_address;                  // mm_interconnect_0:UART_SERIAL_COM_s1_address -> UART_SERIAL_COM:address
	wire         mm_interconnect_0_uart_serial_com_s1_read;                     // mm_interconnect_0:UART_SERIAL_COM_s1_read -> UART_SERIAL_COM:read_n
	wire         mm_interconnect_0_uart_serial_com_s1_begintransfer;            // mm_interconnect_0:UART_SERIAL_COM_s1_begintransfer -> UART_SERIAL_COM:begintransfer
	wire         mm_interconnect_0_uart_serial_com_s1_write;                    // mm_interconnect_0:UART_SERIAL_COM_s1_write -> UART_SERIAL_COM:write_n
	wire  [15:0] mm_interconnect_0_uart_serial_com_s1_writedata;                // mm_interconnect_0:UART_SERIAL_COM_s1_writedata -> UART_SERIAL_COM:writedata
	wire         mm_interconnect_0_gpi0_butn_s1_chipselect;                     // mm_interconnect_0:GPI0_BUTN_s1_chipselect -> GPI0_BUTN:chipselect
	wire  [31:0] mm_interconnect_0_gpi0_butn_s1_readdata;                       // GPI0_BUTN:readdata -> mm_interconnect_0:GPI0_BUTN_s1_readdata
	wire   [1:0] mm_interconnect_0_gpi0_butn_s1_address;                        // mm_interconnect_0:GPI0_BUTN_s1_address -> GPI0_BUTN:address
	wire         mm_interconnect_0_gpi0_butn_s1_write;                          // mm_interconnect_0:GPI0_BUTN_s1_write -> GPI0_BUTN:write_n
	wire  [31:0] mm_interconnect_0_gpi0_butn_s1_writedata;                      // mm_interconnect_0:GPI0_BUTN_s1_writedata -> GPI0_BUTN:writedata
	wire         mm_interconnect_0_gpi1_dipsw_s1_chipselect;                    // mm_interconnect_0:GPI1_DIPSW_s1_chipselect -> GPI1_DIPSW:chipselect
	wire  [31:0] mm_interconnect_0_gpi1_dipsw_s1_readdata;                      // GPI1_DIPSW:readdata -> mm_interconnect_0:GPI1_DIPSW_s1_readdata
	wire   [1:0] mm_interconnect_0_gpi1_dipsw_s1_address;                       // mm_interconnect_0:GPI1_DIPSW_s1_address -> GPI1_DIPSW:address
	wire         mm_interconnect_0_gpi1_dipsw_s1_write;                         // mm_interconnect_0:GPI1_DIPSW_s1_write -> GPI1_DIPSW:write_n
	wire  [31:0] mm_interconnect_0_gpi1_dipsw_s1_writedata;                     // mm_interconnect_0:GPI1_DIPSW_s1_writedata -> GPI1_DIPSW:writedata
	wire         mm_interconnect_0_gpo2_ledg_s1_chipselect;                     // mm_interconnect_0:GPO2_LEDG_s1_chipselect -> GPO2_LEDG:chipselect
	wire  [31:0] mm_interconnect_0_gpo2_ledg_s1_readdata;                       // GPO2_LEDG:readdata -> mm_interconnect_0:GPO2_LEDG_s1_readdata
	wire   [2:0] mm_interconnect_0_gpo2_ledg_s1_address;                        // mm_interconnect_0:GPO2_LEDG_s1_address -> GPO2_LEDG:address
	wire         mm_interconnect_0_gpo2_ledg_s1_write;                          // mm_interconnect_0:GPO2_LEDG_s1_write -> GPO2_LEDG:write_n
	wire  [31:0] mm_interconnect_0_gpo2_ledg_s1_writedata;                      // mm_interconnect_0:GPO2_LEDG_s1_writedata -> GPO2_LEDG:writedata
	wire         mm_interconnect_0_onchip_progmem_s2_chipselect;                // mm_interconnect_0:ONCHIP_PROGMEM_s2_chipselect -> ONCHIP_PROGMEM:chipselect2
	wire  [31:0] mm_interconnect_0_onchip_progmem_s2_readdata;                  // ONCHIP_PROGMEM:readdata2 -> mm_interconnect_0:ONCHIP_PROGMEM_s2_readdata
	wire  [13:0] mm_interconnect_0_onchip_progmem_s2_address;                   // mm_interconnect_0:ONCHIP_PROGMEM_s2_address -> ONCHIP_PROGMEM:address2
	wire   [3:0] mm_interconnect_0_onchip_progmem_s2_byteenable;                // mm_interconnect_0:ONCHIP_PROGMEM_s2_byteenable -> ONCHIP_PROGMEM:byteenable2
	wire         mm_interconnect_0_onchip_progmem_s2_write;                     // mm_interconnect_0:ONCHIP_PROGMEM_s2_write -> ONCHIP_PROGMEM:write2
	wire  [31:0] mm_interconnect_0_onchip_progmem_s2_writedata;                 // mm_interconnect_0:ONCHIP_PROGMEM_s2_writedata -> ONCHIP_PROGMEM:writedata2
	wire         mm_interconnect_0_onchip_progmem_s2_clken;                     // mm_interconnect_0:ONCHIP_PROGMEM_s2_clken -> ONCHIP_PROGMEM:clken2
	wire  [31:0] mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdata;         // NIOSV_M_CPU:timer_sw_agent_readdata -> mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_readdata
	wire         mm_interconnect_0_niosv_m_cpu_timer_sw_agent_waitrequest;      // NIOSV_M_CPU:timer_sw_agent_waitrequest -> mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_waitrequest
	wire   [5:0] mm_interconnect_0_niosv_m_cpu_timer_sw_agent_address;          // mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_address -> NIOSV_M_CPU:timer_sw_agent_address
	wire         mm_interconnect_0_niosv_m_cpu_timer_sw_agent_read;             // mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_read -> NIOSV_M_CPU:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_niosv_m_cpu_timer_sw_agent_byteenable;       // mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_byteenable -> NIOSV_M_CPU:timer_sw_agent_byteenable
	wire         mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdatavalid;    // NIOSV_M_CPU:timer_sw_agent_readdatavalid -> mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_niosv_m_cpu_timer_sw_agent_write;            // mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_write -> NIOSV_M_CPU:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_niosv_m_cpu_timer_sw_agent_writedata;        // mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_writedata -> NIOSV_M_CPU:timer_sw_agent_writedata
	wire         mm_interconnect_0_onchip_progmem_s1_chipselect;                // mm_interconnect_0:ONCHIP_PROGMEM_s1_chipselect -> ONCHIP_PROGMEM:chipselect
	wire  [31:0] mm_interconnect_0_onchip_progmem_s1_readdata;                  // ONCHIP_PROGMEM:readdata -> mm_interconnect_0:ONCHIP_PROGMEM_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_progmem_s1_address;                   // mm_interconnect_0:ONCHIP_PROGMEM_s1_address -> ONCHIP_PROGMEM:address
	wire   [3:0] mm_interconnect_0_onchip_progmem_s1_byteenable;                // mm_interconnect_0:ONCHIP_PROGMEM_s1_byteenable -> ONCHIP_PROGMEM:byteenable
	wire         mm_interconnect_0_onchip_progmem_s1_write;                     // mm_interconnect_0:ONCHIP_PROGMEM_s1_write -> ONCHIP_PROGMEM:write
	wire  [31:0] mm_interconnect_0_onchip_progmem_s1_writedata;                 // mm_interconnect_0:ONCHIP_PROGMEM_s1_writedata -> ONCHIP_PROGMEM:writedata
	wire         mm_interconnect_0_onchip_progmem_s1_clken;                     // mm_interconnect_0:ONCHIP_PROGMEM_s1_clken -> ONCHIP_PROGMEM:clken
	wire         irq_mapper_receiver0_irq;                                      // JTAG_UART_DBG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                      // UART_SERIAL_COM:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                      // GPI0_BUTN:irq -> irq_mapper:receiver2_irq
	wire  [15:0] niosv_m_cpu_platform_irq_rx_irq;                               // irq_mapper:sender_irq -> NIOSV_M_CPU:platform_irq_rx_irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [GPI0_BUTN:reset_n, GPI1_DIPSW:reset_n, GPO2_LEDG:reset_n, JTAG_UART_DBG:rst_n, NIOSV_M_CPU:reset_reset, ONCHIP_PROGMEM:reset, SOC_SYSID:reset_n, UART_SERIAL_COM:reset_n, irq_mapper:reset, mm_interconnect_0:NIOSV_M_CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                            // rst_controller:reset_req -> [ONCHIP_PROGMEM:reset_req, rst_translator:reset_req_in]

	NIOSV_SOC_GPI0_BUTN gpi0_butn (
		.clk        (in_clock_bridge_in_clk_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_gpi0_butn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpi0_butn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpi0_butn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpi0_butn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpi0_butn_s1_readdata),   //                    .readdata
		.in_port    (gpi0_butn_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                   //                 irq.irq
	);

	NIOSV_SOC_GPI1_DIPSW gpi1_dipsw (
		.clk        (in_clock_bridge_in_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_gpi1_dipsw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpi1_dipsw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpi1_dipsw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpi1_dipsw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpi1_dipsw_s1_readdata),   //                    .readdata
		.in_port    (gpi1_dipsw_external_connection_export)       // external_connection.export
	);

	NIOSV_SOC_GPO2_LEDG gpo2_ledg (
		.clk        (in_clock_bridge_in_clk_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_gpo2_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpo2_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpo2_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpo2_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpo2_ledg_s1_readdata),   //                    .readdata
		.out_port   (gpo2_ledg_external_connection_export)       // external_connection.export
	);

	NIOSV_SOC_JTAG_UART_DBG jtag_uart_dbg (
		.clk            (in_clock_bridge_in_clk_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                               //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                       //               irq.irq
	);

	NIOSV_SOC_NIOSV_M_CPU niosv_m_cpu (
		.clk                          (in_clock_bridge_in_clk_clk),                                 //                 clk.clk
		.reset_reset                  (rst_controller_reset_out_reset),                             //               reset.reset
		.platform_irq_rx_irq          (niosv_m_cpu_platform_irq_rx_irq),                            //     platform_irq_rx.irq
		.timer_sw_agent_write         (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_write),         //      timer_sw_agent.write
		.timer_sw_agent_writedata     (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_writedata),     //                    .writedata
		.timer_sw_agent_byteenable    (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_byteenable),    //                    .byteenable
		.timer_sw_agent_address       (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_address),       //                    .address
		.timer_sw_agent_read          (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_read),          //                    .read
		.timer_sw_agent_readdata      (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdata),      //                    .readdata
		.timer_sw_agent_readdatavalid (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdatavalid), //                    .readdatavalid
		.timer_sw_agent_waitrequest   (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_waitrequest),   //                    .waitrequest
		.instruction_manager_awaddr   (niosv_m_cpu_instruction_manager_awaddr),                     // instruction_manager.awaddr
		.instruction_manager_awprot   (niosv_m_cpu_instruction_manager_awprot),                     //                    .awprot
		.instruction_manager_awvalid  (niosv_m_cpu_instruction_manager_awvalid),                    //                    .awvalid
		.instruction_manager_awready  (niosv_m_cpu_instruction_manager_awready),                    //                    .awready
		.instruction_manager_wdata    (niosv_m_cpu_instruction_manager_wdata),                      //                    .wdata
		.instruction_manager_wstrb    (niosv_m_cpu_instruction_manager_wstrb),                      //                    .wstrb
		.instruction_manager_wvalid   (niosv_m_cpu_instruction_manager_wvalid),                     //                    .wvalid
		.instruction_manager_wready   (niosv_m_cpu_instruction_manager_wready),                     //                    .wready
		.instruction_manager_bresp    (niosv_m_cpu_instruction_manager_bresp),                      //                    .bresp
		.instruction_manager_bvalid   (niosv_m_cpu_instruction_manager_bvalid),                     //                    .bvalid
		.instruction_manager_bready   (niosv_m_cpu_instruction_manager_bready),                     //                    .bready
		.instruction_manager_araddr   (niosv_m_cpu_instruction_manager_araddr),                     //                    .araddr
		.instruction_manager_arprot   (niosv_m_cpu_instruction_manager_arprot),                     //                    .arprot
		.instruction_manager_arvalid  (niosv_m_cpu_instruction_manager_arvalid),                    //                    .arvalid
		.instruction_manager_arready  (niosv_m_cpu_instruction_manager_arready),                    //                    .arready
		.instruction_manager_rdata    (niosv_m_cpu_instruction_manager_rdata),                      //                    .rdata
		.instruction_manager_rresp    (niosv_m_cpu_instruction_manager_rresp),                      //                    .rresp
		.instruction_manager_rvalid   (niosv_m_cpu_instruction_manager_rvalid),                     //                    .rvalid
		.instruction_manager_rready   (niosv_m_cpu_instruction_manager_rready),                     //                    .rready
		.data_manager_awaddr          (niosv_m_cpu_data_manager_awaddr),                            //        data_manager.awaddr
		.data_manager_awprot          (niosv_m_cpu_data_manager_awprot),                            //                    .awprot
		.data_manager_awvalid         (niosv_m_cpu_data_manager_awvalid),                           //                    .awvalid
		.data_manager_awready         (niosv_m_cpu_data_manager_awready),                           //                    .awready
		.data_manager_wdata           (niosv_m_cpu_data_manager_wdata),                             //                    .wdata
		.data_manager_wstrb           (niosv_m_cpu_data_manager_wstrb),                             //                    .wstrb
		.data_manager_wvalid          (niosv_m_cpu_data_manager_wvalid),                            //                    .wvalid
		.data_manager_wready          (niosv_m_cpu_data_manager_wready),                            //                    .wready
		.data_manager_bresp           (niosv_m_cpu_data_manager_bresp),                             //                    .bresp
		.data_manager_bvalid          (niosv_m_cpu_data_manager_bvalid),                            //                    .bvalid
		.data_manager_bready          (niosv_m_cpu_data_manager_bready),                            //                    .bready
		.data_manager_araddr          (niosv_m_cpu_data_manager_araddr),                            //                    .araddr
		.data_manager_arprot          (niosv_m_cpu_data_manager_arprot),                            //                    .arprot
		.data_manager_arvalid         (niosv_m_cpu_data_manager_arvalid),                           //                    .arvalid
		.data_manager_arready         (niosv_m_cpu_data_manager_arready),                           //                    .arready
		.data_manager_rdata           (niosv_m_cpu_data_manager_rdata),                             //                    .rdata
		.data_manager_rresp           (niosv_m_cpu_data_manager_rresp),                             //                    .rresp
		.data_manager_rvalid          (niosv_m_cpu_data_manager_rvalid),                            //                    .rvalid
		.data_manager_rready          (niosv_m_cpu_data_manager_rready),                            //                    .rready
		.dm_agent_write               (mm_interconnect_0_niosv_m_cpu_dm_agent_write),               //            dm_agent.write
		.dm_agent_writedata           (mm_interconnect_0_niosv_m_cpu_dm_agent_writedata),           //                    .writedata
		.dm_agent_address             (mm_interconnect_0_niosv_m_cpu_dm_agent_address),             //                    .address
		.dm_agent_read                (mm_interconnect_0_niosv_m_cpu_dm_agent_read),                //                    .read
		.dm_agent_readdata            (mm_interconnect_0_niosv_m_cpu_dm_agent_readdata),            //                    .readdata
		.dm_agent_readdatavalid       (mm_interconnect_0_niosv_m_cpu_dm_agent_readdatavalid),       //                    .readdatavalid
		.dm_agent_waitrequest         (mm_interconnect_0_niosv_m_cpu_dm_agent_waitrequest),         //                    .waitrequest
		.cpu_ecc_status_ecc_status    (),                                                           //      cpu_ecc_status.ecc_status
		.cpu_ecc_status_ecc_source    ()                                                            //                    .ecc_source
	);

	NIOSV_SOC_ONCHIP_PROGMEM onchip_progmem (
		.address     (mm_interconnect_0_onchip_progmem_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_progmem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_progmem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_progmem_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_progmem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_progmem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_progmem_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_onchip_progmem_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_progmem_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_progmem_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_progmem_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_progmem_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_progmem_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_progmem_s2_byteenable), //       .byteenable
		.clk         (in_clock_bridge_in_clk_clk),                     //   clk1.clk
		.reset       (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze      (1'b0)                                            // (terminated)
	);

	NIOSV_SOC_SOC_SYSID soc_sysid (
		.clock    (in_clock_bridge_in_clk_clk),                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                    //         reset.reset_n
		.readdata (mm_interconnect_0_soc_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_soc_sysid_control_slave_address)   //              .address
	);

	NIOSV_SOC_UART_SERIAL_COM uart_serial_com (
		.clk           (in_clock_bridge_in_clk_clk),                         //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address       (mm_interconnect_0_uart_serial_com_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_serial_com_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_serial_com_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_serial_com_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_serial_com_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_serial_com_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_serial_com_s1_readdata),      //                    .readdata
		.rxd           (uart_serial_com_external_connection_rxd),            // external_connection.export
		.txd           (uart_serial_com_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver1_irq)                            //                 irq.irq
	);

	NIOSV_SOC_mm_interconnect_0 mm_interconnect_0 (
		.NIOSV_M_CPU_data_manager_awaddr               (niosv_m_cpu_data_manager_awaddr),                               //                NIOSV_M_CPU_data_manager.awaddr
		.NIOSV_M_CPU_data_manager_awprot               (niosv_m_cpu_data_manager_awprot),                               //                                        .awprot
		.NIOSV_M_CPU_data_manager_awvalid              (niosv_m_cpu_data_manager_awvalid),                              //                                        .awvalid
		.NIOSV_M_CPU_data_manager_awready              (niosv_m_cpu_data_manager_awready),                              //                                        .awready
		.NIOSV_M_CPU_data_manager_wdata                (niosv_m_cpu_data_manager_wdata),                                //                                        .wdata
		.NIOSV_M_CPU_data_manager_wstrb                (niosv_m_cpu_data_manager_wstrb),                                //                                        .wstrb
		.NIOSV_M_CPU_data_manager_wvalid               (niosv_m_cpu_data_manager_wvalid),                               //                                        .wvalid
		.NIOSV_M_CPU_data_manager_wready               (niosv_m_cpu_data_manager_wready),                               //                                        .wready
		.NIOSV_M_CPU_data_manager_bresp                (niosv_m_cpu_data_manager_bresp),                                //                                        .bresp
		.NIOSV_M_CPU_data_manager_bvalid               (niosv_m_cpu_data_manager_bvalid),                               //                                        .bvalid
		.NIOSV_M_CPU_data_manager_bready               (niosv_m_cpu_data_manager_bready),                               //                                        .bready
		.NIOSV_M_CPU_data_manager_araddr               (niosv_m_cpu_data_manager_araddr),                               //                                        .araddr
		.NIOSV_M_CPU_data_manager_arprot               (niosv_m_cpu_data_manager_arprot),                               //                                        .arprot
		.NIOSV_M_CPU_data_manager_arvalid              (niosv_m_cpu_data_manager_arvalid),                              //                                        .arvalid
		.NIOSV_M_CPU_data_manager_arready              (niosv_m_cpu_data_manager_arready),                              //                                        .arready
		.NIOSV_M_CPU_data_manager_rdata                (niosv_m_cpu_data_manager_rdata),                                //                                        .rdata
		.NIOSV_M_CPU_data_manager_rresp                (niosv_m_cpu_data_manager_rresp),                                //                                        .rresp
		.NIOSV_M_CPU_data_manager_rvalid               (niosv_m_cpu_data_manager_rvalid),                               //                                        .rvalid
		.NIOSV_M_CPU_data_manager_rready               (niosv_m_cpu_data_manager_rready),                               //                                        .rready
		.NIOSV_M_CPU_instruction_manager_awaddr        (niosv_m_cpu_instruction_manager_awaddr),                        //         NIOSV_M_CPU_instruction_manager.awaddr
		.NIOSV_M_CPU_instruction_manager_awprot        (niosv_m_cpu_instruction_manager_awprot),                        //                                        .awprot
		.NIOSV_M_CPU_instruction_manager_awvalid       (niosv_m_cpu_instruction_manager_awvalid),                       //                                        .awvalid
		.NIOSV_M_CPU_instruction_manager_awready       (niosv_m_cpu_instruction_manager_awready),                       //                                        .awready
		.NIOSV_M_CPU_instruction_manager_wdata         (niosv_m_cpu_instruction_manager_wdata),                         //                                        .wdata
		.NIOSV_M_CPU_instruction_manager_wstrb         (niosv_m_cpu_instruction_manager_wstrb),                         //                                        .wstrb
		.NIOSV_M_CPU_instruction_manager_wvalid        (niosv_m_cpu_instruction_manager_wvalid),                        //                                        .wvalid
		.NIOSV_M_CPU_instruction_manager_wready        (niosv_m_cpu_instruction_manager_wready),                        //                                        .wready
		.NIOSV_M_CPU_instruction_manager_bresp         (niosv_m_cpu_instruction_manager_bresp),                         //                                        .bresp
		.NIOSV_M_CPU_instruction_manager_bvalid        (niosv_m_cpu_instruction_manager_bvalid),                        //                                        .bvalid
		.NIOSV_M_CPU_instruction_manager_bready        (niosv_m_cpu_instruction_manager_bready),                        //                                        .bready
		.NIOSV_M_CPU_instruction_manager_araddr        (niosv_m_cpu_instruction_manager_araddr),                        //                                        .araddr
		.NIOSV_M_CPU_instruction_manager_arprot        (niosv_m_cpu_instruction_manager_arprot),                        //                                        .arprot
		.NIOSV_M_CPU_instruction_manager_arvalid       (niosv_m_cpu_instruction_manager_arvalid),                       //                                        .arvalid
		.NIOSV_M_CPU_instruction_manager_arready       (niosv_m_cpu_instruction_manager_arready),                       //                                        .arready
		.NIOSV_M_CPU_instruction_manager_rdata         (niosv_m_cpu_instruction_manager_rdata),                         //                                        .rdata
		.NIOSV_M_CPU_instruction_manager_rresp         (niosv_m_cpu_instruction_manager_rresp),                         //                                        .rresp
		.NIOSV_M_CPU_instruction_manager_rvalid        (niosv_m_cpu_instruction_manager_rvalid),                        //                                        .rvalid
		.NIOSV_M_CPU_instruction_manager_rready        (niosv_m_cpu_instruction_manager_rready),                        //                                        .rready
		.IN_CLOCK_BRIDGE_out_clk_clk                   (in_clock_bridge_in_clk_clk),                                    //                 IN_CLOCK_BRIDGE_out_clk.clk
		.NIOSV_M_CPU_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // NIOSV_M_CPU_reset_reset_bridge_in_reset.reset
		.GPI0_BUTN_s1_address                          (mm_interconnect_0_gpi0_butn_s1_address),                        //                            GPI0_BUTN_s1.address
		.GPI0_BUTN_s1_write                            (mm_interconnect_0_gpi0_butn_s1_write),                          //                                        .write
		.GPI0_BUTN_s1_readdata                         (mm_interconnect_0_gpi0_butn_s1_readdata),                       //                                        .readdata
		.GPI0_BUTN_s1_writedata                        (mm_interconnect_0_gpi0_butn_s1_writedata),                      //                                        .writedata
		.GPI0_BUTN_s1_chipselect                       (mm_interconnect_0_gpi0_butn_s1_chipselect),                     //                                        .chipselect
		.GPI1_DIPSW_s1_address                         (mm_interconnect_0_gpi1_dipsw_s1_address),                       //                           GPI1_DIPSW_s1.address
		.GPI1_DIPSW_s1_write                           (mm_interconnect_0_gpi1_dipsw_s1_write),                         //                                        .write
		.GPI1_DIPSW_s1_readdata                        (mm_interconnect_0_gpi1_dipsw_s1_readdata),                      //                                        .readdata
		.GPI1_DIPSW_s1_writedata                       (mm_interconnect_0_gpi1_dipsw_s1_writedata),                     //                                        .writedata
		.GPI1_DIPSW_s1_chipselect                      (mm_interconnect_0_gpi1_dipsw_s1_chipselect),                    //                                        .chipselect
		.GPO2_LEDG_s1_address                          (mm_interconnect_0_gpo2_ledg_s1_address),                        //                            GPO2_LEDG_s1.address
		.GPO2_LEDG_s1_write                            (mm_interconnect_0_gpo2_ledg_s1_write),                          //                                        .write
		.GPO2_LEDG_s1_readdata                         (mm_interconnect_0_gpo2_ledg_s1_readdata),                       //                                        .readdata
		.GPO2_LEDG_s1_writedata                        (mm_interconnect_0_gpo2_ledg_s1_writedata),                      //                                        .writedata
		.GPO2_LEDG_s1_chipselect                       (mm_interconnect_0_gpo2_ledg_s1_chipselect),                     //                                        .chipselect
		.JTAG_UART_DBG_avalon_jtag_slave_address       (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_address),     //         JTAG_UART_DBG_avalon_jtag_slave.address
		.JTAG_UART_DBG_avalon_jtag_slave_write         (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_write),       //                                        .write
		.JTAG_UART_DBG_avalon_jtag_slave_read          (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_read),        //                                        .read
		.JTAG_UART_DBG_avalon_jtag_slave_readdata      (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_readdata),    //                                        .readdata
		.JTAG_UART_DBG_avalon_jtag_slave_writedata     (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_writedata),   //                                        .writedata
		.JTAG_UART_DBG_avalon_jtag_slave_waitrequest   (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.JTAG_UART_DBG_avalon_jtag_slave_chipselect    (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.NIOSV_M_CPU_dm_agent_address                  (mm_interconnect_0_niosv_m_cpu_dm_agent_address),                //                    NIOSV_M_CPU_dm_agent.address
		.NIOSV_M_CPU_dm_agent_write                    (mm_interconnect_0_niosv_m_cpu_dm_agent_write),                  //                                        .write
		.NIOSV_M_CPU_dm_agent_read                     (mm_interconnect_0_niosv_m_cpu_dm_agent_read),                   //                                        .read
		.NIOSV_M_CPU_dm_agent_readdata                 (mm_interconnect_0_niosv_m_cpu_dm_agent_readdata),               //                                        .readdata
		.NIOSV_M_CPU_dm_agent_writedata                (mm_interconnect_0_niosv_m_cpu_dm_agent_writedata),              //                                        .writedata
		.NIOSV_M_CPU_dm_agent_readdatavalid            (mm_interconnect_0_niosv_m_cpu_dm_agent_readdatavalid),          //                                        .readdatavalid
		.NIOSV_M_CPU_dm_agent_waitrequest              (mm_interconnect_0_niosv_m_cpu_dm_agent_waitrequest),            //                                        .waitrequest
		.NIOSV_M_CPU_timer_sw_agent_address            (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_address),          //              NIOSV_M_CPU_timer_sw_agent.address
		.NIOSV_M_CPU_timer_sw_agent_write              (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_write),            //                                        .write
		.NIOSV_M_CPU_timer_sw_agent_read               (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_read),             //                                        .read
		.NIOSV_M_CPU_timer_sw_agent_readdata           (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdata),         //                                        .readdata
		.NIOSV_M_CPU_timer_sw_agent_writedata          (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_writedata),        //                                        .writedata
		.NIOSV_M_CPU_timer_sw_agent_byteenable         (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_byteenable),       //                                        .byteenable
		.NIOSV_M_CPU_timer_sw_agent_readdatavalid      (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdatavalid),    //                                        .readdatavalid
		.NIOSV_M_CPU_timer_sw_agent_waitrequest        (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_waitrequest),      //                                        .waitrequest
		.ONCHIP_PROGMEM_s1_address                     (mm_interconnect_0_onchip_progmem_s1_address),                   //                       ONCHIP_PROGMEM_s1.address
		.ONCHIP_PROGMEM_s1_write                       (mm_interconnect_0_onchip_progmem_s1_write),                     //                                        .write
		.ONCHIP_PROGMEM_s1_readdata                    (mm_interconnect_0_onchip_progmem_s1_readdata),                  //                                        .readdata
		.ONCHIP_PROGMEM_s1_writedata                   (mm_interconnect_0_onchip_progmem_s1_writedata),                 //                                        .writedata
		.ONCHIP_PROGMEM_s1_byteenable                  (mm_interconnect_0_onchip_progmem_s1_byteenable),                //                                        .byteenable
		.ONCHIP_PROGMEM_s1_chipselect                  (mm_interconnect_0_onchip_progmem_s1_chipselect),                //                                        .chipselect
		.ONCHIP_PROGMEM_s1_clken                       (mm_interconnect_0_onchip_progmem_s1_clken),                     //                                        .clken
		.ONCHIP_PROGMEM_s2_address                     (mm_interconnect_0_onchip_progmem_s2_address),                   //                       ONCHIP_PROGMEM_s2.address
		.ONCHIP_PROGMEM_s2_write                       (mm_interconnect_0_onchip_progmem_s2_write),                     //                                        .write
		.ONCHIP_PROGMEM_s2_readdata                    (mm_interconnect_0_onchip_progmem_s2_readdata),                  //                                        .readdata
		.ONCHIP_PROGMEM_s2_writedata                   (mm_interconnect_0_onchip_progmem_s2_writedata),                 //                                        .writedata
		.ONCHIP_PROGMEM_s2_byteenable                  (mm_interconnect_0_onchip_progmem_s2_byteenable),                //                                        .byteenable
		.ONCHIP_PROGMEM_s2_chipselect                  (mm_interconnect_0_onchip_progmem_s2_chipselect),                //                                        .chipselect
		.ONCHIP_PROGMEM_s2_clken                       (mm_interconnect_0_onchip_progmem_s2_clken),                     //                                        .clken
		.SOC_SYSID_control_slave_address               (mm_interconnect_0_soc_sysid_control_slave_address),             //                 SOC_SYSID_control_slave.address
		.SOC_SYSID_control_slave_readdata              (mm_interconnect_0_soc_sysid_control_slave_readdata),            //                                        .readdata
		.UART_SERIAL_COM_s1_address                    (mm_interconnect_0_uart_serial_com_s1_address),                  //                      UART_SERIAL_COM_s1.address
		.UART_SERIAL_COM_s1_write                      (mm_interconnect_0_uart_serial_com_s1_write),                    //                                        .write
		.UART_SERIAL_COM_s1_read                       (mm_interconnect_0_uart_serial_com_s1_read),                     //                                        .read
		.UART_SERIAL_COM_s1_readdata                   (mm_interconnect_0_uart_serial_com_s1_readdata),                 //                                        .readdata
		.UART_SERIAL_COM_s1_writedata                  (mm_interconnect_0_uart_serial_com_s1_writedata),                //                                        .writedata
		.UART_SERIAL_COM_s1_begintransfer              (mm_interconnect_0_uart_serial_com_s1_begintransfer),            //                                        .begintransfer
		.UART_SERIAL_COM_s1_chipselect                 (mm_interconnect_0_uart_serial_com_s1_chipselect)                //                                        .chipselect
	);

	NIOSV_SOC_irq_mapper irq_mapper (
		.clk           (in_clock_bridge_in_clk_clk),      //       clk.clk
		.reset         (rst_controller_reset_out_reset),  // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),        // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),        // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),        // receiver2.irq
		.sender_irq    (niosv_m_cpu_platform_irq_rx_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~in_reset_bridge_in_reset_reset_n),  // reset_in0.reset
		.clk            (in_clock_bridge_in_clk_clk),         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
