��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���-ײ`�>��썅��NX�6�h�@.C��(n)�dm���R^%��ĵ0Ț)���dxÐi�"���fk�G��P�7H���,ߗ�ť>�9�'�m/�Z1K�J��<��b$x��fx���'��+��2Ӥ��J��C��y9c�I	(%F����W�qj%{�o�4a�">�����8^�o)9�/g��M���.�e��-z$����Ac保�NM��5�Y +�6�����p��E:Y[��_�xT�I��r>���g�l�������,pS��b���ļb	�R����/��	8�j?��6
���7˳9�Z�v�G
��5k���:�S�ME�XN:�j.3%����5�Pk{��Б_�&��u�m�k�`M�`���p'�f�'�l�l��qaQ݃/���4)Ҫ��1`O����3�Y��[-�
j��g���m笽mbI��`�}}�pk�xyG��)|�wD�������~�RĮ?�*X;�d�KG�;��
�q��d�+K0��5Cz6��AYy%�&Q��<� "�?�$�H���H����P���{"����ZWx[�1�����N�jinԜ���k^��,��5�ղ�o���>_c���$�r$2�J����Pr�T��W~�e�O��<�r���&�t7�?60���?.���I��yP��;���Z�E��Ha�O4�9����=���ˣr
�匑Lg
dwV�(�C�q$ �.�[&��(�=�)��*]߫�HE��Y����f��aqP8`��r�q�Sw���I���(yZ��WOL]�ת�վ��n�5�*:~��9?�$k��~���d�_�t{�_���r��r�� ��M7��I�u��P]�6_߇p��9��cG�������.p���������6�e�t�=��^(����ҋ�ۇ���=]ݤ��ý׋8ƖU�]zͫT�?��ZX��v�#f�mo.���+�\��̰��"�=;#(����Ep�I��w&�J9�R�K��fY>� _"��U�s��]�+�D �����ۚ���������H��q�{�w*�4����/J
�V��%~��#�*'���YҸ4ge��rQw��Y�o���_�t�H�sx�0�b\<���ʹ��؊�T�����[Z=v�t�ʹ���Q���9$�Z���l�_rv?���B��J����F��`g�5�`Tؤ� /�K������3t�:Y��x�֧\��%��F��P�2����,%X�)e���b�g1�����Y�D�RD!���l��O�X�K��zJ6%�C��7�!��3��D^�츷z�Z��%�p�|{(�l����,s���K�{wl4^:/��݊��~�ܛGuҵhDW�����/[���� ��6�i5��I!`����:�n�@����5��	�v�0gw��-:�6aW-�ɏ䇢V�:�U=�	���%#A>ȹ��qr�}0�ۀ=�v�13�Ӗ��(����c�_���a���2��3#��f�$;�?WjU�M1�w��$X��#'K�~V�ƀ���1��8��C���寤7�F��p�S��4�Y�&���,
��e�JU�o�����vcD���͘z(��1Zɿ�*Jֵ(V�T����e�(�f��&վ�z��Q�ܺ ��@Fpa^��<�6CGݏ\\�G�Kwu�:D�������2Oy��){Q9 �3=/}s�cHT�;��	a�T�\(�#�eô��C��GƖ�<��R�7������>��gڿ#��3��̈�;\�e���� W<o�y z��*0�A$(�״�-�mi��QDVq�,��-��V��2#��#���AP�W��IuWN�q�+��~&~�� ������?T:	��K�N_��?��<W!�)'���ƾ�f>W�[����\����&8��B��g�3��މlu�I���Q:]He�R\߉a����U���v]�8sd ��$�@����Df[֜ �u����?�Yq{l��q��t��A����9���}�T��Q�,�=شC��0��~�O8��Ac	���V8�'����%8ᕽ,��͚h��;�cUE*F�
X �]<�?P���#2�yv9,�yj ��Ɛ����&��Ut�\�g����m�	RO����~^��Y	]��~�_վIK���q���-)��>��n�$������=
�v ���5��7��҈��C����-�>�\
>\�:����� �v8(D��­b��Z�o�`q|I7����[��S��}.ǋ�
y�m�:'$������`��� ��@��ٜ�V��WE��v�u������k��;�P+�$� �h�.��ӣ(�!��%'�d�:?��� ��~���9;PX���?���#����7~_&��HY8�D\,���j�M��4����R.a��;��g��ha%�9�|�>���b���s�!M�,�^.��H��������m%����j|<3m�:�2a����S�n����|�-T�deP��z����1�-�������=ձ�y�����/¡��sP����5����I����}����.?��0�1��n��y�[�q0@n і8���<�S[���h�5"�p�$�j���PZ�rÚ�I�l@���ϼZ�fX�� l��<
/�/n�H��l���t�ꆰ'Ƴ��`A<*c~��u�{W�N]�ݙ��a����s��sO|hqb�_�
���P�gih;su�TQ��WP�D]����]��o��$��F�1�@��؀P�GML%Ȍl�n��_�1�3/p�>��^d�f<�7&��WXm��7J�ASɿ]ub��N��!�%��,�I*k��=��m����&,�IMb@9�]�e�E�@f@t�K���ܪm^��F�t�	��^e�o�X�	���O��X0�[f�|�E���W����Ҳ@{�Fr�)�$��C��y�#0âa�n�5�R��%�����G���U>�	K�*�*u�j����w] ����?�ft�'v�
�ܙ��^X��"@^@{�B��D\1�̌������ފM�JW��4,���*�J>�򺞤�ٖ�46��"��qS������) e������1[ڜMn�U�6��eV/�Eb� y��b.���1�E�V���h("�� a��5/�搜N��h�����Z�����$���P=����s�c��?Ҟp���@ĊDX��xM"Y�(3�Fv�N��.�ǡ��e�X7[,4�އ4���\��N���/�a]5��I�W֔���Zl��o�鼡Q�]�,���(pPX�yΥ u�Ss�a��l�N�SA� w�1�g�5�U� ��V#1yh��"���i:�(\^;1%��x��$�#��X��Gg0����wN�r�0���@�o��8��v����T�� wѨ�)rr�oF^�ٶ�:Ƽ��Cd&F�!����38�\�b���;��h�x�0a8
 ��7X��":��~Q/1n�+:�Q�� F� )O��g�$��ؕ4%�s+�b����)2�%�r�^H�+c�%(cJ���AfH��lM��B>vUI�ԒLI)�=-ոF�1�GF����x�K&�A|)J���]R�<�{Vݷ�̗Zt	�ӑ�q 7���YʼǤ�X^Cx�0���s��+��J0P��J@���Wml�̤4��⁔�"���q����o)������h��B*�� ����kK=C�����=B�fj��N���ݽ�˝��5NB�.����&����2���(�c5��ǡ���
ui7xʹ���9�y��y.��bh��t�j�%�/�}d��>8S�)jrl���x���]1R�Xjl!;�(�ךu��e���ұ��VCvP�?E�� �w�����n��`�}'8��yt*���O���?��(���[�۶�!�;-�`������kN��<
u��"8�u�gc��"h�h�S�u�-H��~Tm���n��b1j1;,"#:��/��5��}�Z	h���.؀�v��S1B�]�z;���#���N��B����5<|L���+<n�^W�G[�����T.�ޓ�_/Ƭ��������B��J�@LVu'�CN_'}�!?:���cr��c�^ ����dw�>>K=��hC����rk�o=e���$�lhn��䐭Y��a;����Z�{K�Xk40��M��S�R�̪���
R��qF^���z@^~�G�<�̠�=�v�]/+5�D&�H�kte��wF5��ɰ�{	�/&�֤4�vYB�d���䨥s�L�%�gk9Wp(�ݴ���g�SB��t���$<HB��Jt¦ey�;7O��e������qA�kJ�H����q/`Ј�a�x��c&�d�F�$d��n�/T�$<%���vN� q�l"a��$��.��7;)/"�7�S���zl0�V�_Ç�H&�u��&���q�X�N� xɼ�K{�r�>����m/�j���wۘ8@N.L���{�����vYM��ho�t7H�P���p��������ܱ:�`�{Ct&�Whq1>����r 5$iֳ�} �줠��z�����mHkp��q�ΏSj�h�o��߄N/r�~�:R���Q}2>,�Y}�Q�"6%'�J�����z�0"��rul�*��%	`R��� �r��.-�U~°���t���ֲ�C�d{5�D�d���2RK����|E�S,�|D.�O�]�#uƽ<�}|��էf���I�K���xku(P�I��PS���w4������11[�#>#�Z�y]m_�OM����^��XRd����mѣ*�������S��1UĪ�Y�l���=	�*�]LM�@Ii$�ƍ`��7�+(0�b��  ��,5��m^x�:t�����;��=��`��w<�l"��>�F�հҴ�������٧��b���%�}�V:��t�����5HU?R��g����y��i�Av�$(��wc���Se���I�����V�ƌFܻm��P'�����_x���#1�ez\P�5f��5T��q����d����&���l�pl���j��M�cJa��x/�@�nT�HR����(��A1b����U���O�`s�6�e��B��w"�Np"�����٢���������Y4Մ8k�|����=zˍ�-�b��7i�,��x=D����`>�,��G��N��(>�Z�����[Ŷ��5j��\��=9�[���>�*3�8�Nj��$0ِ]��(W�	N¿-�t���gxlG�dl����� ��Tݷ�ê�ce�@p���\��k6�`�)��w�z��g,�6��I�� �Q���öJj�&�����B�Ƕ|<\�%Cc�Ha]!�`f4d�<͘�׼�E�Tՙ%1��W_�O���N׏+ݍ�����ν��pS哉�0���������l�1�0���Z�/�@�j�Z�y���!�q*�L�)���N�	�|��r�M�y�<Ρ���t}�����*�G�tqܓ���H��\g�2�����&��/L�iaEj��!JC��*ٙ���n�@��ߋlQc%T��vɬ"�`5�xn�����"�����E)�=�QW/�*0i����y0�FQ�TM�?��]e��+��e ��5��2Rn�ESW���*��nw����G��t�AYU&��K�1��v+������ڤKA�=~��z�X��y\�ц`�a��f��k����c�cRGB��y���?z,TMO�㶪�geӅ�KԀ��Y������K?�����~R{ǘ��k{�i�B:m�v�R�ohM��n��A��+v�˴@s:�����§�GI�!�����-�1���o8\N��M�'|z���֝�8:�y�?�ZTY������è��k� j�k�"So�ו��r�H��
��8����]
���[DT�	S��vۮ�r��%���S���a��*$�ajY�3yu�c�uh���t�'ԙ�X)�"c� /uD��������on��hy9�+��w,O�>����� ��_�"���Q��W��{�����)ȅ���W���Ҭ+!k�ۿ�-�g5l����˳�0є�#V��&Uq���>c�,�N6F:?ΨnI��.b�"IO�\:�YcU��^i����D�9<|�Ώ؋)ǃp��yI�'.s
l���َ�	W@��#�������A��r�J��ue\u��v�&+�ꝰΑ(L��y���Z��9�6�iFM�=Y�s䣫n�b�����l]u�p�0<�|���Na�j���1*������G��լ��|�J��l��K������Q���r $����X�������u�ޖ�3����!���#�觥G�{X9`��?�nȱ�SźQ�f'�f�V�Ğ'�Z*O�=��Ҕ և�Xw�F�C@{Dt#dN�ٿ�G�]M)zv�%�a�~Y��@�+��r��a*��(0#��s�@�s�������RbE_a���G���')M�,�;_@ ������=�����>Sw^����ix���OD�B��x�|s�ņ���f��w��緌`ŠP��
r�=������-��������M#�n��vxNo�������b�l�\�O�}�+���_�sN��rp�`a�s�~`��R	��깚�;a3m�	O҈+�����^]F�zK^��$��Q)���"!"��Q�z��8�52�܏̫�4#����Q�K*,���]�C�����������b-s�q6��̴!�|Ns��#S���*��,�����R�N����yV#s+:
�����0�ȿ]�����	��&�H).�E/E����U�țt$��w�#}�Z�T��b�R9��r��_�n�J�|��c�*�a�׹�3�w]B�P޸@�.�Z�߿���^C�H-ɸg}G~7I i�摭=�N<�Z�n��&>eX���A�6nb�H���ղ���l��j�*�_ʄ�3x3ٽd�5!�OF�B��0�(�|�pN�j!�Q�4��C�� Q��X��n�a|Q5��T�O	O��9���Uw����.or.�Z�uF��+=a�p�h�E\=����q�!4���+NuZ4JFs#��'4͟;�2�Fd��ID�6�G_�3ye����a��-��s�ƾ�w��Z{� �fD��542��5D�r��L�y��9<�i,�A��9r���L��3f^z�@%��.Oe�o��p �
l7q�>��P�^z� +�u[�9�Xpuu�4_�'2N8�"����m������o?x[���KZW�B%Sr��Ӏ�W������Aawx�p��h1]f��t-�Խ� χϋa��>əy�m�I�VI'2�@;Y��7}3�	���{#�#�a�(a�b7�V &��s
PX�Ri����̷��MKJgA�c��9�hn��B���	p���H�m�h\I���^�+;��釼H6tk_& ��7�5�&�~IM�Q=�c�d��9�U4KZ�yY������ܜ�
[%��rBĤLԶ�s��#U���=���_������jD���p U}��U?�<�T�?~`ɾ�%������<�����<��ǂA2-�|l�臖v]�S*��b��|��qoђ*�?0��C��$-���0P���ܡ�%* �~�� �`��ο���[��z���2�����[%6���J��\�)�=R���M��vf-7`� iN�ƞ2�QgT]A�*ê��٭�|9!(�Fb������j���.%c˭
����8�xNu.چ�w��[�%q��e�b؛/RB�>t���/.[�鎡�gl�ږ��5e��)t;�@��
�(�+��TpT�*��J$:��KA��`\q ��\�.k.�nقg<�b��AQ�Y��Ŗi�p~�a��=��y�j�¾����܇�;�8SA�������h���)>3�Q5���͐]�i T��a���>�l�gy�����NsL�
$J}Bm�Ԯ\R�H��8��:��b{Hǭ^��O)m��X9_N�g����".<�^�&Գ@�. ��	p�Q�9˾����q��g��ٝ:ؤ������+�m*�Ra!J�����E��h�4Jv����CS�9�E�eK���U��aD�/0k�|���Ď�5���W9+�H0�q�@�γ�-r9�0�7��y/E�������@���ӕ�`�t�
�y�͙�'-w���E|:����K�Ng
�����vӁ?q�ԣ$��jyʷ�9K=ƣV�(;���m������N��L.����NH�RF(�p����`����ų�=�c-���+0C� �.�~�m�w�4f�� ���t!�G�?�7�5�ԑ��͑֝u���n���y}�5&s����	�b����k���#��p@�q|��k�쮨NO�87��v˙K��λ$	�-oNgpD�|�y�ƌ����<|�3���d�ε�H�Z�C�og�0��=��Hr�U�y�Z�@��sF\,Z	qz����4���� $e?8~m �L�u 0�	����]�5�!"�'�<f?ב�����g��h��צ�q�X�q��E�N=��S5�� |w�k��k7�#�*%Q^�߰E<��g?ǂy)��C��/ۧD��nE���LPWus��MlIIe���d��,].��.}C[t��_"�-`@���+OLg��Y�Ǥe�X�uܣ[g0�Qڕ�V���A�eY����H���k��dQ�z��h�TwC(U�d��g�Y@K��;C�ʀ3~��w:j�/n8�5_��e�@�^e�q�f �ۃ,K���"ӱ4�𮼋��2Ӟ���t�\+3&���Q�?�E�m���A� ���%���N���|���4�V�5�(��q��K���lW]P�c-+\��T
h��D�����D��H۬��3���~�a3��#f�!)%�9��ȜȼE8�e-'V�]/�PC*�D���.�~�0F�ؚ��&���[���>��?ɀ���V�����)�'�d�����8B�k#L���{#8<�ق2}V�r;�~�@���-��W�yL9��Ծ��k�R�����C��ōc�ʳ2��/��(�����^t��Q��" m�n�f��0X�����W��N[����5態�%�t��ٹ�A@\��AO�eO�� ��g�2�>@�of�o3�SӺ�Dz���D��+�,	��β;��~�h� ��	��P��HS��"�m�j�4�{�{�T�٭�e��$}���:���#� ��$�k���u�����`�a���}%7�B�D-��o9d���sT\���/^~��wT�B��uQ(���?���������d���|Ʀ�$]�q_\�����\`�:�˱[)^�	v�P%1ߵ@` 	Cj����<Zn@v�/a9�h��sP�99���c�ds2��D�ED��z�{�� ~O�����'��HԂ�o���{ϟ|�Qq�{lA}�'��wT�ޔE�I�k����.�b9I̓�ë��&�l�7�>˃�8�_bJ���|ua�����@��c�b�t}���]�A��VR�U"��r�2~�g����?���
�"���"D'6{�����z$��c���������!Dw�V԰!`9���Q+�g���:P���u�$H�g�h�1�Q~�$ծ˭}�H�Ќ��Ut`��5��\���������/.Zxn��©'֘��57}��5��B ����t�T�%ӭ{J��P��^��"�����#���Cbfp�)�{��BPk��n#�ͽ����+��$|^r����m�د	�
���7�Wm�c0E�VE5��&}��R�D���P+]�$�|�7������h�Ψ@$)�D{PZ�M���늕�k��zw�*�>�e�-���C�H�'a0�YGؙO"�ǳL/f��d��\kG�0P��h$0`�ߕ�=��V����b���[T� 6K�Z�����@|�2�n9��]���+�ؕ�X���;��W�NEв]� \G���.�i�4�~M�'K�ZE�F���	������,gs��K�F�^7C���8�c�2�H��c�ٿ��D@S��	�~���C�,�L^��:g����8]1=��*6����MU