��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a�����/�	v�+����@ɧ-3�����Iz�t�܀Le'H>	6"�U{��9�bEɤ6-�!�V��s� ���m�|����~μn���}�iԹ*VC�4���m7���-� �7�o�d�0wUQ�z:F��:�����wq9NI�|�'����b�C��Ӥ�I��Cz��,�7Xmf7D��3Y?&L3�?j��h��o�dƛ�0��H��A�H'Fp؍TCP����W��p�/MBq��� ��,�NG��Ӣ��:�6K9R�d��Hf��o ���]��0/���Q�'�FȨ)��V7Ⱥ̀;"ݰ����g�,I=��^?i�S�@)�h��P��4��+���'� )|<v��$�i,�)����Tw����~A,�i��Z�lput�?>��U���T�)"R���F��	&j�M7����G��~�?B��\���jj2�#WK;������!���]_�ڇ������`gF ��jΥd���HrG�
ܶ��?xX�,0�Ֆ�'MĻ?���} ��X�@�o��l$F,�)�IOqV\ݨԯ2y�Nȫ�D�>^�XE���VQaCp������a�~7��Zbu���/�cB�h�3Y��Yw����VO �/C+2kT*J!8-��?\�N���X(�?c	S���5R��P��m�R�´����ʚ�&e0�G�x�d��&�ZcfN8YjQ�!��K�iW1�s ��¶�pT�dв�t,�&��䫓d�Z�`v`���V�qFE�T��E�·\��� ���`��1�`�b a�D�.��;�����VBsC�"4��:gƔ�Qт�I"UR"`��҂/��T͠� q@_)���A�Dh��qG���U,<�	h��v�0y[FzJRH��,�Z��kā| ����Kp�/q��B�N1Kd��}r�U:�Cb~�P3�R��o�h�+!Ӓgb�S�0�ήSg� �^V�}r���T,�V�t&��y'��Մ��T�l�ڡڻ�H2���<���ˁ��2Clw	�����?�p��Fw�9R/�LY4��Ʀ��z�M����`I�9�:�ELn����Q��ۥ����J�Q���r�[�S�S���M��<N*#��5�}+_��M��ؚ��|�5\H��VPe��ِ�x��@/L���53q~n�W��̲���ȕo�`Ьd=c(�j��f'��X1,u.0���Ö� �t\��$��"����x-���KA�ԥ�1fvȠ�$t�l��[���TJX^p�>,����fh�n�K(ӡ2󧦣����,
��E3��j"�ԓ��r���)F>FTF�~��D9��}y֒��j�#��E���ax4d��p <�b��=��f�:����lvk��DwЀ7����J,�%@ۥ�L��b yl>�>>��>�D��>��N�^= #j��*�7�ZA�h!�z`�	��@K��/�ܓ'R0���z����$0��.���F�Jj��hRk�mYQr��&!�ƨ@9Y4�AQ3<�+�*YPx�N�>ðM��:^��]	a�Q ??O��G$��dl�pt���x���z��ڊe��Rkh�Y���EA��\M�Eh��$`��|�'"�R�ݒ2����ma{(tRW�Q�����]a-c�F��7������)O�]ʢHK�~� ͱ��0evĜ���je[SK����aQ�s�[:U���H�CAw���/��}��	����l�:��bM�l�������5?�<
D����c �r�V������N�o��l�%R�U��8,z�wZ����>�9����2�خ���$��|�)�8��i��zx�!�xB+A�o����Wq(	k%w�(Ռ���i��P*`�O�KFֶ����H�1[r4n���C��o�E(��6&ʕ�@f���Z>%�BJG�@����d�+��J�_��m��
�=�>����Q�i���X�9(sM�'�H�n�C������f���6�n�C3���V�Y9��\��܉l�EUܑ�I��b�ęm�ǌ����h��.J������qm8{��4��'Vʇ�*�Nh0�KaF!�-ha~�:3�����@p�cD��l�Pl׾9a�ML� $����@k`l.f�<�'頖�誑|@�ճ;�G&~(�N����[�C��;���"���[��"��Ω%�i޶�'�_M�}}Z�����"���V��`"I�)C�0��x0q��`�DӲ�c����k�ǐ�@�&�&�[���q˰T/��)�e�)�x)��U_h-�{�M�`�Z+�]wp0C��Q��,lwj��
� ���e/���3�Dc�NS��ȣ�n�,؅g�_�)��i���<�Hob޺��}�N|v%��hQ�LU�/��NѤܞ�X��Xe=�Εb�h�ڕް�a��mG�[g�&�7[Τ�7$nW����Z�	��lw�TTk�n(�c3���ʛ�'��p���^Қ־��T�� ��ڣS�C�rps8���YJSNڿ��7d+���_��v��A���zc*T��ER�� ����$���vvJ���c��h�y@T�����}ȴׄ�qD�a��mT=;)@+��j#z5ku�ep� 
a����>�u��p(l��wYSH$�;�ʗNy��7G�(�Ʒ�=�3Oa��m���Z0kji9��='RAH��i=s!r6�9����;q���F�\����d#�#	'A'����a��A7��jF��!�#�YM%|�F����<gf?=p ���Z(n���W�B.��ܿ�5:���v�B�S�N8�7ء
m]&-����-�6����m�;T$j�������o
5�|b�y���U��>&'���S�]t�dE��Vp�
?l�E���}OzI�@Hwz^��/q}�_V�<B�^��؁Ejxj�{����%���-��si��/��g�����1��JB�޼�qd�n@1Mc@�����%Ǽ��1}����*�Nq�4_,�ﳤ�(��K'�b�c�E�<6�ĝ���b�I�r&P/f������b|���h-|��7&�f��H,�\�;��l�0Z蒍��E����%�P�lo��GO���>�^o�(Fa��TU���D�*9�Ej��h�"5��GQ�5�n22�ʞ�lz�~�}����˳b��9.�aw/ ��&�;�ڌ��Mx�xq� ��S��E/��d����e��ǐ�1Jl��)^4N��5?=9�kN	�҂���g}�Zo���e�Wi�E�����\�˟�Cs_p���Q��~��hq�1�.���
��^|�h+�;MZUz���4o�J)I_���YO��x���� �˃ �=�|�z
���At�b�תި"�з3M|�J�%�u-�d-�/�!4ю&5�{�@�y?o�U�Dȃc]�{�~�'�ߺ���AG$����+<C3�;��B��8W�{�EE&��XQ
3NS�B��UE�sw��h4�Ig/(]";���˅��4����8�����g����@
z2�l��I����`St�=pZ���>{���`K�L�,&��lƉ�����]�2E�σ����3�ϯ��o|'K�zF��O^Q�C��4��������@$��&,j�r��	�1��3�8�%IW�,�ȡ-/lN����K+k�4��01�I������5�"�4USv�\fn����qߘ���N��L;�h�&K)i[���筱vzk]x�#t�R���������DԈ�c�F$A���1��+�6L��hb��ƨ�q�Z����"�� ,\U��2>b`Ӎ%8�����
��1܊����G{1�-��-�'k6=p�Y�^?E*�JYH�4�%x������A�=8�;��sx ���N��������|�+��y�qNr��u#S(��mk�?�����"`U'o<��$Yn��cIBx�{_����3���������Z$Y������O{��a�Fρ+��^���B�<�Y0�Y�N�P�����6���9�^`�ߚ��|Y�2�8�!����Ŝ�o���x�W��H�k����ܹ�j��YS�4e����-�~��/'o[���/ta�_���0:Y��Z��� z��\tͲ?-���d2�d� A$��Φ��FO���s+R���v%��Р�1�܌�Cƛ�bb�q�`c�U�,߶ڵ�M�6����x��W^��@o�ʉa(�ކԶq =��0��9�gv��{�/D���ϩ��gs��}���<�'�E��A�A��#��<
��"���bB�pK����_�A,S26F�iy�wޒ��{�ǯ�)DҠ�ԅ�6�)�>�:Y����[�^��]y.��{�odQb4�m��䭗,�鈊=Ds-�y�K���T��%H�p}�`xE�\�������Ɉ`(xr���s����m:ֺN��U��
j�*e����� Q0�N�u�ԣ����V���\K�s��!~T}�yE�����춄AX�w��G ��{�"�(�{�32kn1����2F��
����{㏎�!B��M���s5�:J�V�F�З�qd���C��g~��Z��1!����|V���Po�x�+�E��J�f���,��^��[��O%����h\��GqZF���3/���f*0��`�2F�~G��QmXUs�1��._9�0�U�HN�����ni��,]߹���.�e�u��1yH�rv2�dIZw�J�J5�q���g�Y>�ZR��slG�Q^ɿ�����6��l��\kV>q�{����\><��А���E��4J ))&L�E!xገO7Z�!��a21/���d�����(n��=3q ~	/��v]�IV�,N�A7!Wf=5�|��I�!�wz�0&zQ
��k��9l�H$����R�mq�_��r@���q�� ��/��`����na8ohu8hwʾ*P:D���>��|�cs_�x��Z�ư���3v��U�n�c�S����\=�:�o�QTO�}�h�mYs�n<�+*�ј��V=]C*ou�:�(/�>^����ZL N���C�[ZKm�:��p��s��T��Pi�N�0�ƞ�L��d?�i>O�l�~�X����=�=����a�[��O�٠�C�(�S��_6Y?�����Pͣ�0P�t� (Ft$/��gC��c�`�4�8�)s��I�M�((��)��4C?yt�w_>1����߮C`�wCǱ��D��On�hdY{lT�H�C����t���yH�\��3"�ϔ�u�,3�ǫK�Og< �s�.����J�_�
�s�?�B01�G);� ���S���;a\!��N��d�6�����x�#n��L;��ʦ~�_3���%T��hhn�� хxPIO�q�*��Ѕޯ��'28z�s�l�wk�ADi�f�s�~��֝@�nϷ��9����E�`x�[���Z�q���$*E73���(���1,O�S1�~L�,�R&ϗzG2�K\ۍ ��m%�U�?�VVޙ7YE_N�X:���ɒ��x��C����D�i��w`^۬��R�pk�r�u��.TS
��M��ï������R�-�hĆ	��|�*� ^���#ޱ*0(�T&�Hq�<u�⾦�кm}�.V�.V>n� �WAUu��P��t/- f��{��Y�O�i�I>~��y�42�3�E���YJ�x����
�.,cqS��g˕]��V�Dk#��ڛ�����[3�::e
�I:�+������o#�D�YY�:�oz�����F�~�څ[����i�����:VG﫮5̯
Tb7�M|tV����K����֤P�9oѤ���\1���Cq��@Pq)H]ţ�T��Qa�S������֛.�W��Ϫ?�$��M��M�7���z�m�~k���^�A��vR|���km%�AC�7礦�]f{=-�J������v��C���RU
�kÅ�86���;�B�����]���?}��GBa�>`
-� }����dk�;y�RR24rS�9����zG_��HM������� ���VT�z:x�7Y��$V&=Po}$�ø�x���r��`Q�yt2��{�J�|�ޒ�c�.�����rF��j��-NL$�q�Ֆ}�� 3YT�Vx��#T�q�l,3�a��.�{�͸Y��Ҥ>�j�sAj��Qk�M�/�P�Vc��2�a��~kB������8l(#�ʔu���3ʌh���o�l��������������EJ�����m+�U�+���7�j`^��������)��sn���׊><r(P�+NŸ	�_�T��Xi�_�u��5>.�����8 g@�ӆ�C���0T� �8bXR��$8R1_��'JpL����1��u+S��F�~��~��2N��ɍ5��G�	���b��H�[��y&
k�|�N�}�%�jף.����ï������G>!x��c ����h��p�)�_�m��V�Q���i�蠮�P�D뤂6P��F�l>����HK*�U{ժw��� ����(X ً�-�S3@3<ｸ����UH�Y&S{��f��0j��E"7�}������
�W(AIY۴D��?5��b�Kb���Z�jsbVp�1�Z��X/��j���O�O�I�x��������0z�FNl�ZT��S�d܇\i�$v���	t��2�+���"����)�ZM.�WCCNY��a���PK*ȗ�n2#�R�odj���o2�i����L�fT����'���
�ƕsً�YmN��5�e��#����w�fidy�S ���oȴ��n���a]����s�s��>����)��2s�FK��N	V�r�gŝ�OO�H��#x���E��  �?ݨ߭-׶aݮ�3>9�.e�[x���`��ڳ�72�\]�,�z"A����л���)�oQ�*�&��@<��Nx2��V��&)�'�P�"G-ns1��Bf$^���s�!�ОS��R�#`�םv�L���D^��Zi��:2�H������^����w��ꚯ�9�	�� ֍@ǲ�m����{r,4�*�L�/T��>��g7p`�9т��vx��*p��S�ty���C~�p`��3���Ts�Mp�S$�� �u�vQ����(5�	�9�˳ۦ�N�B���¿_�[� $Xc/�M'z�j)��f�с�5�Ҽ��CT(����P��@lћ�����V7�sC��f���Џ���	Kwho!)�~��V�zP�����.��4 u%Y��*�]�6IW���Pf�VcD�v��۲����w��s��~��OW�k?r�[Q_��&����@�{DC�*�5�.�&�[�6˰\/��q�[�z����#�
l��%�@|�;�Ŭ�J� �@|�����63��[M]�S�j���H�M6�c�=m�
+��"����񏨅����i��3w`��}QY :Ho����CP�=�_WC�f��۶�ơz��/\�w���i�丁�=H͔~���+�#O��g���ٝ�UD_��c��v�؉�v��u����>\{x�&���>�A�6}�Uk�>�����5��U�r	NKR[xӼOI���M���]c�!T\�6���s�LB���?qYkZ99�.#9?�WdV:Xz�;��	~txCR��)���Q��?|�P����r��Q��Z��s�\x�X'{��%��Ws�d�(ǋ������Q%u�ݚ�xAnC��kD�B��s(��y�8����̭�d��m-N��,;�9(���W���z�S̂]� �~=���Lg 6'��4��ٺ�J���ql��?��(N,�Q�Uso���4$��2.a�Z�<��;;�ϯ�QZ����iuZ5�g|�!H�<��&���O�:B ��g}Z�O�O���5�\(��hve���*�� kr!�e�r�{�����B^^V)�P����}Y������k����~7����y���8(Ax���?��C�"я�6D Pp���О��WL+4��Eݤ8�. �ځߣA�����o,Ӷ)�2]�<+38�s2
�mTc��^���#��<,�t4���mp�zM�����*�ӭo"�a���"x�E�w�6���i5��p�*�GwY�����Ki�����c�H�×p莩���cMG�U��Syo���9ԑrw_y@�ʛ�C�r����4�}�w�h����Z�ժ�I܉���Ft5�[�Z�~3��-�P�����[3c~q�3��9��.=z!ݱs6�S#9��(��{C�v��f�����`�E���Natی�U�����D�p��I#
��9TԫH:X�e5�E�u2\\Y�~yz�)���Y��o����}���z5����!f�}9���Aei�KKkmψݺc.8�s�[�/�X�֟�DWIF�"udG��ϊԻ�t`ݣ��`���6@��A��C�c�^PB��H�FQ
�	ɿ5�K3�|�Y�;o*������?H�, �z�H����<�3`
����eK`B����Մ9���(sG�8�&���a}�e���ӝ�E*T��:�Mi"�=Kt}���R����&_��۬��̫Ȇ�#��q��j]��%z&�=�[.@'
']Ol�]�_�7���\wHխh$}��Mt��y��ڀJbwuڱ��[5�dH�{{�n�Z�� ^}Z���O����H�E�3F�����~�W��� ���ҹgA��3�?��%�z�:�[f�_�h���'�>\����`��K]�9�,���+��=�&b� � +��WiS����Xh���?�!�`K��;�9��==`��\gc>u�2�����w4�P��ڽY&���Cװ� �G�j���nf^�0ASn��*�V�������E[�����>�n��s0��QJ��"&�`���/�a�5�I��w"2��%��L=Oۆ�B�K8�����v��ez����uΉ��0l���)[�Cv���e2K�S��:g�'`HDˈ��њ���#(�"�x��'���.0�Ww�$��3�y��?Qu�V}5d�;�� �^[ ����ʞ�0Zs(0��Am��D�.���@��/k;��wA�r���C<<�m��g��E�� ��)�!3�a�-�3�F�e��O�F~��RUw}Iy2�?b��m6�,�M�ـ���%RC塮�=@8���!�N*]�V�'ߖ/�А���;���!��O� �
�/��}X�U����?J4%%pp	�:�?{�<r$64�(��m�D�U�,g��C��D��"$��?��+�=6S1aa�PEZTz ��!�7GA��]+����Fy�
�}�N���kܚ	hK�Ae�� }�H�xo�y�x[ g��\�r�A�hQ�9�=�Ǥ`c������?���2�MV��O54�� �!�����V�P]�(�b��sK�P�����nx�G���A�dPS��,���1���h�;��i4�&�Q8
�ܒ���?X�P5[#�_����|1��~� �[�ȧm�M#��&�6�[���tOa�6r�j�����
�z.*����s�}��K�<g���|GmL�"�x=fҩ�5RH��OU2kȆy$l�Ո���B��UM��<F�������q>�Yi��J�^�_�Re�p�����
`.u��c6R}��NjH|	�� ��/�;.�y��H���"�٧�:��s�g	-<�vsb%vyr*�`��d�������I]�7o���nG��S��ވ�-���G�], ���F<���5�.�v%k��-�q҅�]�����J�1u��[Ɯ(�:3���Y�k�4n��Q?@#xݣ>*�7RMۏ鑧I�%g�����(#\q�D�����%5y
����`�+���&��I��2�Q���ʏs��_�0���{�����i-n:��'57��5�V���\��zC���s8u1,,�Rב�lUX�^�ǟ5�cbhf��ĸJ�(�ScZ���Fξ�cC� _��"x��ڲA��Go�8e��95��w��)��K����>F��ײ�m\����2�^B�b��	�іm�����r�Zߌ��)O\Άw���-��;c2��/qX�%5�N2�"ggi��C��W��[pym���є�I�h �6n��R���ޯ�,<����Me-����.V��2���zԈ��y����(�N�DY���a���X�#�X�<��`n�M7�O����	}��۲yp��k6:f"��q}$+�B��G�Q���E�옎���cձ����w[ӥ�S*;��J���2�zƭ!���u�c�����3��n(Y�;ÉK#�q���aoY�w9ܥ�m�Li$h��������@4u	4�J���r����l�"�@�e@0�ڊ�ښ�E��^����.:�}�
�Y�N�?<��4,
3��[�ȥ��@	EgTE�\6�T{���r��5֔'�@x�+T
#,�J�,�#�ߢ'F	6v��#6��P��,Zm���c#�����0��?b*̝�uC|vT���YA$�\�8�*TY�E/d���bk�I�3��;d���������d��Y�J��@�M�]�^M�~��B �fI9���R�����q��R0�ꪇ���?$���Dںe
�%5�������=���S��yQ���b}6�ݿt/�K"ɷ[JUi@�tk�ba�XK0���w4��,�~vs�Q �c'?�B�N��y!�nw��2�պt�`�]6J���óM����϶�Zo�J�i�����`��d.��x䤚U'��P�#�J�*&����֤�N� 貺��U�
t�3{V�ڽp���T
�H�K�'�]�I6G]$"�S�w�zh��t-���PV.��5Q�����m.g�"f�e���<�}�wO�@��c�z*��a���%~�3���.��fso�r�}L�)��Y�u�m3�;�A;?��@���©��}��'�&A��
�E���Bf@C��mܘe�,����o�^����/y����H)���XS��ݯ�"�ݔ�T�n�O.���t�*����e#�/�G-Hh]�-P�����7A���\:�=�����RO��T��-Pk���ɗK/�t��m9����Yw���&�A�[;�(�E4~��ш�QBF���x�ضA�5�ȳ��1��a.3[!��Np���ط�F���f'������j%{>�+���e���
.dH���bD�ꅓzU�"�s�T/hi���ܖW�ӭ�������X<���K��+�N��Ւid��W)X:B�*��.�9�=Rae8�c�qct�r��5��I�}>Z��(QD>�V��!��4+�ټF��)V�,Ua
�3���ua.ő��rd���L�2�2��g��V`E+�����J�t�orzz&8ic�P���~G9�X�A(�,{�f�J����Go���U���_h��x�U�D!����Dua����H\���(�]w������b1����:V\����J��r9�T�8;�\��;����)O�\a����ֶ]�еk��G|�r΋qR<�u�Q���q��7���ؖ@��Px'=��!��
�/Fi�m�5�1M����ؔ��@;�Y���9���~zH���R��t��D���	3��<������7�A����vl��r�sl"�i>��F,㗎N<4ʩH��&
	�-�NS�_��پ��Ƨ*�A?�4�/�K�Vfs+�y��~Rpu��0�ʅ���T�]Q��%&�8o��q�t�֪��9��O[��	K8|���s�ah�Z���8�����F��O��`�~Aj7-�Aͤ����a�]���(I��f���J�6E�������$fּѷ�%�+e~�\	�?�4,�ai��hY�5�� h�0��1�8d�ʐ��+p +��(m �d<�<���j�E�33������B�Ą�J��P��2���R痹iǔ>t]������J#�앗�p�[���@��F��G��ȶmo�\ ��Zwm��]e|z��ݠq�ey8kȵ-+�E|�/�m�ZO�q���r30�g6�/����n2���/�8����}d8�(����w�M��i���k���$���ߴ����K�:�~��^�4�<���O��,ԫ�ݞ���Ę�rjS��n��F\ǥp-�3A�������XǸx�Dq�����
+���������
Ik�h��fH������t�I�qp��!�4n�
�4Ȧc�����lpdܻ�,�Y�6�]��4E#V�ɓI����&u0�z����� ����ɍ/0�t:�"Y�y�r�i�R�w8J��	�����ڀ:0Y�u�����`��V����"��:�AŮ?�<1�.% [��2� 2�b�YI]t�;�W�T�fZ ����&�,BL��mT7����JG���4��.W/�*�bL�&b����i�4�b�H��
kv"
��fN��}> L����ٖK�0�_�-��~�}:/1�QЀʈ�:I�ͮ��%)S����b���/�=�z�i\��
���#X�;���0V;��犌��M4�Ђ�+��\�=d�H��B̂W����2hz���φ#��)}i����6��Gʗ6��~�V��\�lR_>g�T�5/y�������癮S�Uް}o����tent��-��,X���f̙E�e5ÀJtNrh��||������}�>f�}�m<:�����I&�e��
��Q��2cm��YxB��=����'&eʖ����������J&uT����xr�g�W��j�`jkĘ�`��������&����z�mu2�닒���y�$�t������`I��鰓�{�k���>!�͒;�zdx�ID}F�c�T�u��l��O:G�`)(�����00��I��v�i�_���W
O]x��_��Q>�m����p���X��V�A+�sj��m'ZA�{C�8�e�����IU���@�j�!�O�{.v�9���!3M�ܺFd�艭�U���޵��	�E�h& A-U͡:�4���������� i�A0�^ɠ�`�:�o��� C�UL�����K�K7�{�7�YiW(��%m�)����f��)����0z|��
��])�"�1k��P�V��$A���1̴Rr�+ xS��*��	� Y�9��K7t�<�-9�����ޅ���9��"����Q�H�s-Uy�"�9�5�LZ���&��-6�L�H�����u�/q�V��7X�Q7��<*�?k<��b�r�S���\q0�K�;շ�LXۇ_�^�b�"�ޔ�Mk�}y�j��1��3�Q:m��HytƄO�{�a�
7sRIH���[؀4�ba��'���R֋7HQ4-iO>$Sت,ʫ�Pa��4"�D��@w��Io�xg�T]�4���4ם�g��i"��d��9T�iԘ�	;=`2J��pXg�Ѐ���ƴNK����V�L	��C`��>3��_~�z�4�v���-��)ŋ
N�`�����+�����e(Ɏ�zQ� �?G#��e���"f����8�I��ub@X�.�0o�6T�����MI�w��		��.9��#����|�������X^���N�Tsnp��W�吁�?#����.����Ͻ�Y ��):RUݖy	� ��L�0���{�F�S[�+Vq��X�n�DFz������3*�~=��6�z�ߪ��}�[q\�:f�@H���9�������ǧ��I��J�(df�c!��u��\&5�ƚ� H�c��	K�wJ�� U��	�
5>�r��p�\5�e=n�5�&N��"��=`-E9�y����A.�/<b���!$�r�T�Yj}lO��̯?*E�w����F"4S� ���݆Ds��D߶t֟5�����߳H��3Aȑ;���䠑�8�[\4�Z�kq��� �jUXB���ű���+(�d��Z�a�{�oŇ�:9�p�����s�5�6�tؗR��7ވ�0og3pw`~VW{�;]{Z�ީl����M�ɖ;*�KEb<T�3��������O{5����@�+���������G���2hb�[9�"��v2�O�t���c=g��$�.Cm�5��z�A����!�#
��~������{�]�!{ 4a� >�T�E+B�����-��d6Wb�ⷛ[oi���WZ��&��q�;�Y��R�$]�Y���]�Fs�=S&!R�/�EƩkg�'�'��mw���bi�Q �����s��cf����En�|�ٰ�3��.�a�1���w�^	_��ԉ�����|?��7�W�3G�)���/ r�r��g��g��`ml���4�\8�&L��Ы����B�&gAT���3KKg�5xG�|�k!u�D�(�57�Ee�vX`r!ܨ|�O%�
�lGc��X9Di�p*��)v���%ΰ7+�HL��?�-l⟖@'���v�xڥ�����0��6s�b�3�l7XO�[�\�c(hҮ/ބTب3����W��b�g����ȕH�́[��,�$w�H���S��}���,���p����ת�Q8|[C�󆮲]�C�3�5�*�y9�ڧ�3�ʇe��,и�u���Jt D�ĩ�J �۱�fq"ǋ�첓�Wi���r+S?d.��繉���`ь/�D���}x�)@�ѺO�5K��b4b�qvn&܂�։��޺�Vfm~�#i���n!�m{|��l��8ӃZZ�X�Q[p3b8��\���&rL⫎�K��$��.�%THd�[�gp8�T�n�u�&]uMU|dL!m
"�W�Re�����[�M�d��l;&�@J?k�od?粍h���ƞ� ҷ;�0�������v5ͭ��SE��%v�'����(��{�*ߍ�g�ҥ�"����H�1.Ƚ^�;��24���[>+~�JFq�#(��+�Q##��#~�.?�6��f�,�Տ��&)�[�x��?��o��`�b�+�Ĥp����L�l�������N��%�Zw���C?�׳=E�=_��`� �ߣ��}{=g���h����"��4'�#a)&�5�Y3��tľ� =Q�c))���V�0#�\ޗ�+���VFM�|�U��8R>�*�3�C�uń�� �����n���|�x*Z�&��n�tֈz�
A��잮y�hca&U���ro�ka���M�W9F��}�*�g�|�7T�2�M�  �&_P�'��p-}uݭ� �oQףGZ�Nr���\�D���U��C��R�0f�������۽�� e\x�Qq�`�o#%�CE[J���b翰)�qa6���ǡ�6�I�RG%J4̉gF�|��?%��@Ak<��S�H	Y��I���8�~�
��X+a�_=�s9:�/)(
� ȿv������|>S/�?�N|�ܣ1��鑴ԍ�i��X>."�<Q�ܽq����;7�Vx�g���dd���Ɯ��|�����8�`\��Ii�3m6�-!��.W��N�G�:X�v����8>8�ܨH�.Yg��5�@��S��T���՛�?WtV���|t�^�V�b�gcd}�G����ٻ��7�ݒb�t>�)թ����-t�<��PK��3�/�a�}5���Y�e�y'|�j��vf�>w(��C�F�t�-����&`6����j�C({�'mش�i�f�v�lf[+��K��>��.[s)1<c,�F"嶷F��6��������J^晐Dr��h]10��HΣ��m���DM��Gቖ�%�QYPJ�� ��%�W֚ʛ9�X����x��F������V�^E�#9C��uU2�s\�ďOu��S�|ob��܆Ǥ��_�LH���a�l����\����e
�%�# oV���Ql�O��/��a�����X�"�j�D����osB�o �5�F:��9ґ#�|f�M�d���,s��u\��m!^�G�þ��{R�ua�g�e �Ԝ�#����m�0�f����AC�N�ބ���ߣz��&`N���� R�n�qF7$dWI{���j�5��V�-(p��n�xq'�엱�����Qd�5|N���w�\����F���{m/�ΘM�);K�w��:���:����N�� 8�פw`�����Rk}f#�n���h�ǐ�[c/���Ik���sY�����큝��l�w{0���e����ua��m Rg�<$H�)��=	jWb�gG�R�b�������Qva�@�]�Y��꧚�!h�n8(�̩"z<��Q/H��&0[�e�He���"��f�iO��؉˹��v7o���b�1�ޤ���[n��ڔ*�O��N(%��JP�+@[1��l�+_��eɷu��b.�ћ���1�ڦ��k\/_�[����1�{�H&D���ˬ�dG6,򟋜9"5����'�d��*<���Y�Ӄ�&ANc�˹Jى����ו�}_S ]21ԅj��;��?�����-a���CE�X zP�Hڻ�4���⺹D�s!D�(���"[�ڞ���@5$�x|>�?��W�
oMȴ9���\G�N���9b������OiE�%\9�&����3��:�s����&?���ɵ��D�mO땼�Y'�[��*�s�?�7�/
vFeZ䟚�"G����|�v��%��G�O����h��k@8}U��݀[�IW��Y$=y	�3/>a�^%?�������,�q
�vM��'��xM�_ �'�s�{Kz�Rڇ2�0��.�&�*�u�X�A���� �W7�;y�J�j��&}&ūX�O�W6AvmmiL+�#O=�M�;.f�5BWzp�e��0�Ȁ�&~|kcx`BT.U�4���?��#�ݥ
�.ރp�lq���`���P��n�P�����
L����0:kri&Tـ���"�`N�(E��W�Λ��E�R,łH�-1EZ*L�Ӄ�l��\z�p#V��76�%��F��ϓHo�&�6Ä&}-*����	���ﱐ"iH��#�}a�ֳ���?7GY	Ր
 E��|e���0X���@{�M�FЃ)��;mcՙnjV �R��u��Ӷ"1_5`���Ȃ��<� l{@3��2�*3n��N)��>4��*�{��>�z���a�ug�K�~rx�'�nL���n��{����高���[<�"3�,�1Z%ӽ��{=��FGX�7c[A�i��qi��5<�d�a�q�([��H4�l
M�Oy�k���-��YHס���g/��_�x��`���k��Ą3��!تe`�t"��m��֍j2M��c������U�ܜ�-K=�V\:nG��o�r�K�P^����X�E,�T��u�;��Pւt�r��6P��Av��եH3���K��h�Xֲ���9��X��@.E�ӹA����"��;��ٝoQ=5����T��X�6x.Fy�Ujۓ�y�t�š��+nV�Zݹ,��ՆeJ_������LQx��P��?�Q������,ޕ�#&1!�q��b�P�Sָ�ゝ,�KAt�)�P� �4�:�X�s.��S_w��d�z��� Zn�OxC�� ���ԟ;�9w�&��^߂s"��9K�|q���D#@*���EkǙ�o��˼e�B4��G7��r30���3�@��V�O�T�=����ś��+�:2ˆ�[�8����.�5=����v�h;đ�.-n��n��)�5�f���:��������Pֿ˄���vZ�@چh+k:���m/ݳ��w���W`V��1��ܘ��u�5u=���:y�Ȏ��jpѡ� ��~�u}[f�-�1����`�씽���[�[��*	���G���,�ӶS=���3с�.�&oj?qo� �?� ��V�S3K�E�[���B�@��)蝫g
��(�<MɧR�����~�y�ɜ���B�W~������z{�GM�7�1?7�� �F䄳S�8H('�3�V�P�I띥0*�z�_�M�yW%¹���ݸ{t�H�V�#v�#�>����q����$B��3��oO�̅$��75�� e2���taL���o�S���)�8y~ۂ+���]k����|�441��X�Hʙ����yc�B�%M	�u@�Q�g+��T��uB���NК��
��P��Mj�5�h�u�w�k^Wv���/k�� ��1��T^�M���QI6|��C��}ӯD-�(i;�*M�I��]L�M�=�iX~�O�xa� �G�Gŵ���a�P4�))�N7@�7�&|gψn�u�}+I+fӦa2ϰ^���g78��p&9��M��k�V�j X��i��U�|؇s�:���uF{Y��m��E�I�}�=Y�]:��<�|�z�����Z�o`��_s!�dU�S��!�㓚ڹ�R��T�D��q�r�7������z�ޑ�״�x�l���	�M�p����<��ISwܭM�H�]���x�{��,f�_l�-��",$G��z�.T0!ͅ�{3�"����P��FA��^xrh�
ۗ�W]��.�`T�8Z�B|S0��>	��cN�myHU2�P�|�qe��[\������ť��4	'��R�o�h,hN"�z3N�"g�H5���*O���Y����9'�����̕�<�?�{��]�;�W�*?,p�ּ�Np}.��(&;!/����_o\�+@"2��]��u�k[w� �5@,�
r@�{!C��P���(�W�YPs3'���ȯp���o߮B�]����A�p�י=�\��}���,w�QMp,��/��ˠ�m�{pE��8��5 �	�C�CD~%���4��'Y����_�� 8�ɀ�-g|�W�O���˘�6���H��Vuݝ4��o����H�Y���?Ig�&���A��f�'2�=����f�IT�Fr�9�|-��G��E)��iK����7A�ۑ�pT�
�p�X��`�T�M�ͻ%$3�%��_��3��jm��S��H^I�tZeת+ ��*�n/�kS�t�� $������TBkH���}]����48���M)@�^6l����f���zڠ���#��iEH}�]���'L����0��p]��8	}��L�g�<` �������D����&Q�er<	�KѰ�(9���3���K�z����$��@����'�:c�L*�U%Ԇϧ䃠܊J���r�)S Y�,�Obq�;�������H2����1����MD_LdCw�a��ᅐ�xN�4���:>Hbb�%E3m�E��bg�D���� �Y�?�t\a�UX��"�w.��X	[�X��Ԫ=2�Ǩc@�x2��1�s�� ;5�y�=y*3A����C����{���nY��q7��&7��a�����֙+�+�q��R�_��ƒ��MZ��f���va'�P��9?CM#��aX�����۳{���DMS0�R��j[�D*F�ms��OE{�o�W?p�Qj2�g��2�p��F�S����Xے0�|��f�𡺐��H9�Xn��u|Հ��`�(�x�U��Ż�ˊ�s҉�����8+�K뷤(f�e�̖����}O�6ϣ�w���h�0�]�m@"$�	���/E(�T��:.�oWl�$���L<Pgz�3zZuJЊ(���d��$�9���F��#0x*>���f��n�I�Nf��,�*�UȒ9�� ;���%��Z��&:k7�z�W���g?��O1?�� j����H5EI��ؾf��C�����i��� OH�u����l��I �4r�j�9J��1�7�<�|=�Vu{9b_ � !��LV+K�dF����X����\��#@�sd�SDm�o9���ԃH">�X�
�?3�]_�F����q�J��X�����x�2ؓ���q�F�C�~�R��2w	6��;�$!q ��h<�T��w�aB1��Ƀř�J�.�%��u��}�ͦQ߿{6I�b��E��$U�X!9�~8邶@{������I�V��ޔ��t,cvD��~�y/��+B'H�K-��0��B?��y7�J�R�(�$4����ښto0�g?�c<�F:��p�F�8�#��y�����Y�ҵ0�m�_�I�\Im�2��r��3:�D��Ѽ�mk��>��,eF�N����w�p�l���X�q���vYi�3�2ʃ�dU�F"���P]I�{AY��G�[V��V�B�������^ ���	���Zqd�����o��B4�?r��kʲ�0���]-�g��S2��D�H�6M�'���KI�R�u�;����c��~A�C�;�N�xB�,���%|���ʧL	��p�� ��?���P�F�,���ӻ�V��?B�/�l/�
�0V�GWm��y����;�4���=��^�a�s�T֠���>��K���+�c�H̒W���v�~!gvc�ȋξV�2i��;̜�ܥU�,E�s6�O�Ba��X����;;��/���a��oN3������d.3�{ѻ]);���C��"��'f�hyF�7�I������5���տ�eg��'�uPL�+��E0�_9��(����{�����_&�ϲ�h�^]�����z���]|)J�}�R쬊���	UU���e8�4m�yTJ��N0��uE���p�*��/��VEɺRU���?mL���V��s��t a�0�8���3"V5�v���k���u緁�9{ �0{��,ϑJc `8����8v�4>�d1�X��$���B���0�)�jG�)a��QW��{ZM�]�Z�^ݑ��v���b���>��Y-�\XtW\�YZG�G�B!Ȱ4���
�W7�V
����{���sڊ��*�aX�����t���z�s�it����D}{��,Ȟ�K/2:��^''
��>���cel��O��SZ���9I�{�^�q��pJd�,��X�� ���j�~;M�Z>Y^��pꖘ0��)|4[7_�&�h�5�|H�n���]�R�_GY3Q���_����}#�L��T���z��� �&��jl{�.�6�Aa���t)5�EJ��eV�ޝ�7%q��45�-���L/r$h�m2F���ܕ�@�\�=lດD�Z,2B�=�P�i���s�rZi���Q걧7�`6�r���_%���J�&�ܭ��B�`� }����b��6VN�����<��1=�;���.�Q�qh�<�p0=)z���`'SP�+�Jn!y��Z�A�Z@�~L��4��IX��ϓ���`0��F;�R� QV��p쇦�-�u�M�~�hT�u���#(�'3������Y�Wˊ� /lf���fA� V���'�*[��6b���o��W�Ѻ�HLopY.4A�2o�Tv��3�?��y��˗!�&,�<����򫱄��$� �������{�x�,́�����{��_��`�}?Z���a��:
@.\�f�Z%Z�~M��J0I��1�����Uph�:�K��k��(��|�
�?� �KW��T�_ 	d*�1�=\>�k�+O�A^�p�s��~E>���B�*ۅ�<�����!&(n����m-�ԥ+��,:�`k禮hd�{Kw(:��)W��AH��v�"	��[i7G��ȷ��4�3�|��7v�����hY�<�]E,��7{D5W�DX��7*I���_�z�i���gT������a��<"���A�8���Y�� �~�3��$�v�5Đ0�^E�4�e�{�⠯�
�=��&BPO'ZBR%Z��u�C���)�x6@����c����L\}�yO��	��D�DB���sαyJgY��8ȝ�}ÎM���5V�� ~�Bu�V�ؔ�f�"�,�� ��*��H���<�6�]0<�}�P�Il*<_��[qנǁ��;s=`'�%^���t�u5�����JK��.0Q�n�Do�ͼ��q ���RټN���po�]�y�+pn69.��!�j��41+)2U�	GX�}�C��q^����X$/l��<ۖ�ݡ�8Ttv�ދ`STN"�Z&�	<�+��zW�"G6�f�$gB4����~��<�\�D���Ǟ�z�~��h��R�rZ�V45(ph�z���g#R�����<�3���|<4�	����=˰Cݯ�I��:؝���i�,l���-�y���/�ui�,��<~��e��i��lr�������Y��s�F�Lx
-[��#xN��0��:j��e��#�>���{���Y�����E]�U6���7�$�C�׷��.�;��XH�<U�bT~����H����x}h��8��d �J�6�� mX�dR2�QmѢ}�S1����,dE	�� "@?��(��%[|��U���'
�*��@˺< 6�g^X����=s��9�[W��jj�r��"�d��1�|��M�e,�
I�6�5:3O���S���%s*���~����q]ݿ�-h��hP�����o1�P6�6s!�����KK�i�4�JW����*��EO&N"��c �5�U����	�*�f9��U��h:�&���v\�v�%ŸF�{ �C���L̽
���*�`�)�^����5(��T��-qn�상0�%E��˫Qf�x�G������Q��������tzw-O.�����4 ��|��ŵ�n��/zz��3e���vF�z5�t���tl84\�d�q�����3�	�����������בfN���5~+�H���j��ܮ[J|��c�8Wc��9~F���x��0*-!m3�c����y;4��|ҷ!k��"�Dں�y`)s��T�/�Y��c:5�����舣���TϏ #s�&�þ��6b�R���ҮX���7"7�}x8�<?����&Z�o>Aj>�-Eu�֗�C0�EJf��N���Q��^�m|yyS��; �4�ݜ��HZ�,�T���X���v�ՃC��?u&H;�&���X������;;O�фl��ް���f|1�x�{�Zb?��d|���þx����e�,20�4�p�<rEP���Oa�҉��%�A0_!:\�5�g��\�^0rl�	�W��O�O��w<���x���7�?	��К�����?��۔�8���%"��p$�l�!�1.q5�D��;&o�J�iR0oGtiPs	������؄&�7`���%�=0��V�e�J@�:S_{�
��F���~'\�%�s��E�KM�V���)�=��V3+ힸ&�_�y���m��b������#��C�Zo�[T�kBL��Qe䜫d����Ćg���1��YI�~�# gr��K�qe�}��O������/�?z��"%a'+)��t��(��t��LZ�<h��X�٨a<��	ptJ�? �נp���$��B W�N����_�,��Ρ8x�����މx����/J�B���)���c�mC-��y��,X�i���,��cQ�X�%K!�uԥ��}�+�H�����l�h&tvu�.�H7#�5���ت�_rU}�/nZ�R{�O8ƹ��]8�	�W��$/�eĥ��@O-����5��m�4��p��z����Uu��c�E>�u��!V!�ﯖ٘�ڗ ����!��
��U^��S�dM2P�K�s�H�O̗?��zJ���Zp��#�f8�z�sq�[��>g����-��SgCv{?�~����4[xS���\�k_�t�J��9��V�}}�a��B��C����$�0M�.{{�{02�!�I����[�G���H�˫揊�.(���mZO)	�h�}F�WA���8/��u���U��F�Q�w41��liKS����*�9sݠ�'��B��my�v�|$O����P��p�Erg�C��D(>��ꡳݭʆo��Y	
x��h �"30EY?t�N�t���B��k��������Y�F�:�oi�;��<�-��*��.^�uM@ a���{���3R�B�6RgEq6����R�<݊��+�/��Y�o<~\(�K�4h ������˲�������'U�W�"g
���%Z�Ĕ��ch��.��hw�
Ș�UJrC��p�S�w,L��t������PDŉ/J��J�s�}{�	�`V�`��}1|��51i�S�K{��Vp��;������E���?B��f���Vb�<�xtq=%�dJ;z^q-<.Ê�`V�oJ~t{��Cg�/Bv؈Kv���zy6hIM5�%&�v7����B`/g��˷dC��<v	� x	���+�O�흕D��6B�Z�N�)�#�M�n��|��ƵBO&�T�}��|#$��k�M�p�<��H�6iߊG��o�Ykpi o�5{��.dV}�T�_�p�Q��W��Å�8���+��c�ht*Q�~N�"�a��Ʈ���p����BV!&��3~6Hf!�-�^r�yp��&��@��p�2)?�^tnܼs �C�.�;
!}��G�V�a����A�eD��ծWE����:��L���U��hG�ċ�p1~g>�dƆYL�c�-b��;W�ɧZ�Y$�BtR6���L�
��čH�H�f:�k50a���#�U�� ��[�2�S�2����$*�H��	�ݱD�+�6/�P{���v�e�c�N���R+垪���oz�3T߾Ju��G X4]G?��t��J]�t̚���(�`�W�<���Xm{�A`8��X�Z��f����/l 9[�<n�F:�NL��~u��3�θ��f���LD@wEdㅗ�V�+ ��Lk�_�'E�Zs%<��@
B��V/*s�O����zXp���	^.ē�hk�|<������n������ʳ�a�����Iy�h�L1c����"i�A��s��C:��1jQ��喲�i-��<>��FB�B/���b�kR^��vj��e��:|'�zT�Vgs9�g��Җ�>�,����=@ L�
{s�3��\��&���TsDC#����dd� ��xo8V���SX����̨��c������M9G�Э�\��p�)hS�!�Ov?Hh��I+�\5����{�GXj���2lb@�vM�9��g���
�?�lW�ޚ6K�X��^%0�ͱ�Tp��t���>/������� ��9GZ>fX~l˥"�8�d�_��^�)�WQ;k3Wʌ�C��`������Z�J�A,��ߧ�F�<D	�
j�s%��T���_�� ���R4��9��/|�[�=	(�ދ��F�9_E��j���t�-P8���bL�6���hf�[.=:�$�	l�Y��Ҍ�����3�V�����K�<P	������Pq�JK�e�����>k2��@�O��ˆ@1��]I�� �{�S=��l��Ā�f��±�\��cd�7��_���	2�Hm��o���Es���!�E�M7*s����x�r~��I�i,�H�}ǩ�V��vVi�&S��B��^�Uhp�[t�ͽ�|�p�k3��/��x�Uh`[,�՗������7Ԟ7\B	&�DEs��{As����(O�=�L d>Ŋ�X�V���M�p�W����S��IS7j�y�βf����R`�������l\�De�Չ!���+�d���2rG33�pmm�'���Бh�P�I�7:m+����j9�?w���Y�A+�8&�+*�������/7�"q%{=ǹ��(���)���A8�aX�Y�`S���!H��Y��84�NP*����� X�ZE��r}](�p�N1a�ۂ�}�:}Z�9�PUi%Ibv���^��߁�Y2�֔���Ƈ-@�9�Ǯ1���c>L]��*��рtP�T�̙j�X��<���0�a���������Y� W3�Ke�}��$y�`�|4S�^��Jj4�H5;��?�]PxllR����c7�4�<���4)U�}X$Y���GSI��ɠ�N+�1H��+E��
�2����%h�5�ݧ�>�bB@3��&Š���=PM�ƙ�O�WvAO��ߓ�mYWܾ*�3�R��A��d�0��B�̣��U�I��j���J'���ȟ�!3B;�M@v��x��fb��Q+��a c���Oz��Y�~Xm��>>a�fRI�tbņ��-�N�-l)]}�Q��|�E1d�y^
�(�JR�S��sy�804eB/�o���ʈ����ڼ�h��;tB`G|��LȒJ���e_٥5��̇��y�D�To4t�F�	s�*�R�}L{�}�����mr�@.��?y9w�hYS8��ʪW
Ђ�\�[�g�č��Qp�4L	�S��kd�(�����R�<Η͛�F'������^�"�^CSG�&z�G, <~�m�3׌4$���N�DN��g'�{Z��$
�q��h��R�g9J�ĳ3��aO���|��,�<R�����tz��3ʧ�Tn���i��>~�L�A ϊ2�F,�Ok|��M8���� ������ֽ����[�P�������ˁ��r�6lFߎ�Ϝ�xs��4���h���45tL �J[�O6h�.]����zg��aIm�c�r&���"�6e�7����J��CO�G�b�e���`�>`�&EFh��MA���6-�K��:��fo�X��n�����C��O�d�I�4�c�ʜ����^�|�a"�7,��!�5&�uu�U��"SU��Fŭ��<#W�3��_���8������[�p��2�c�r��Y!� ���r�l.�.*?����p!����E�/�9�)�6���a<�~~�S?�H�V���Z��p���=�X���!���T�]?��Z'}SS6T�!Ҋ��k�)�|�Yֽ�����czH�y��aq*���s�+��t�$
HT�M��Kcݷ�3l�'�'��� L������������m�;.�.��b�(ɗ`���M.%f7�Z�#ۙ��X`���,�������B�W7a�9_TRp
�9.�]��W�5f�2�(�v�n�vQaC
~�Uf<$�5�Y.;���0DB���3���'G��g�'��)b��\��4�Hn�%���٣rn�a�S�&���c����l��H��T���b��Aߤ��8T%#�����\O(m��7���t�w�H�pmډ2Dg�t@
X�X;cQŹ��"������^Ni���n�3-�+An�@���&j��Q��%h��4���JS��	���s�Fp�������t�R�qĨ���2%����:/�SFk3z���7�oH�u���JF���k��`���M�&����Kj�XR�)�}+�:Or�#�� CY����,�,��ID��P�(rWQ��;�&�c���b��p ��a�|�,���S��h�Ǿ%���-�f/�F��J��A[�h�Q� ����w�ؒ�T�/(8k�̠b���A��� �i��Q��I���#ME��3ۉ��|�7/�<�˹�W�?�O��Dk;'�g�z�kW � ��2~�ܓLq��s��>Xn���x��c#�K/kw>������۬L�-�p�Qm�K������)Q8l��/3�
CO>~�N �2B7�����e`r�z�� y+�2;�4�I����o�;��Q(���q? _{$�7�U�]�Ō|���kԉ�NA�B6�.?�q��jOw�wN��'��������{�W��6
� �s�{�X��2-<v��|��r�*��!+��Eb�!�QX�ex����e�*��KZ#/�����6���,��gn���=�@�>��U;��u
?ݩ�(�pƭ^u9_�~�MU�M���*˸	HնQ|���:�`z@����vs$��e���3�:ʒ��,Yi�m���͞�
��!�R�,J|_����O�R��Q���\�'(���Xg@�����7{[�����GZ(|�_�{�vwG�����)����v��co&���ى9�R�kg%X	���#�XF��.Då���8e��w���3}�9�h��?���[�Y��uY�>�!ვ���r����8wr4��,�$�#`���Ý�q(B���0t����0 h?�we�o8��oq�\��C3��!`���#A��9���vs�z�4�7����Z�g�
j7���e���{F�.@v,�݋��4���UG������ C�B��=W�k��	����ν�jPy�V�_�ɳ����H����/��ZF�-��$̼�<VIl�|V�����>��a�6؇X?������ˍ��i�z��j�Ϯ��p&+<�ǀ��w�j��cR���X<;���֟�}拤Vz�ԣ�/��%a��9i�dխX iLρn2-�� �a� p���G���E�볒�Ĵ����@P��#������%�HR�$0���e�b'���o��GNܩ4(�W�\�r�{#R�c�`PI�6�e
�����u%�2[�ٺ���n!V&4��UL���N s]���6�+�|Yuj�]�òAJ�oȶ��$�j9(�:g�� KڋW"�����eQrg8\�CӶ���-h�'0`?�T��`�H�U5x3���F,�P���$�!��gl�Ԫ�_���b5���d;Ǽ�Bf�G�_h����`j#�!�{���I���IR��ᛕ=(2B�����jҟ�sf�g�T�|�q8�m*��'qԘ�/Ij���X|���5d�(T=+-�w�SA�f�ۇ�9�{c�����s�`�G����xxf_�o/�f�*�̮{���qN3뒯X��b]��d\��U��D<U�����p&�[ ��<U���q���֬�����J�^h��DH�Y���M�?�uWd�(�ڣ*���T6����JE��efS�o���~�An����G���ϻ�it�)�O,��x�[7(� ���	���1���;e5�h�I"�,��(*��X؅�`�O��W[��B�|�x�W���f���j�ٛ���_�H^�5��{�\v!l��7�y�FJ������@��,����������7�][��%�	7�N�*���a�fg�P��h;�����JCۜ�:Hv���Y�{~�T=r'�(4`�}g1c������fn��d:�����UO���O���r1�	D�Ȕ
�g&"y�e;ɹhW���ߨ���}ܨ��I�R^f�|��#2y
E�����%w���!<����T�ѽW雽��о���`|�e�(rk��w0�*t���S
v�}���I��d�7�J�(�9�5�>����{=� zSl��-�ߣ���- 	�3������	��9���q�.�	1��]:��؛tk��J8`x�8&�G��&�Z@G�]�i���j^~�\WqR�DL��t� ���"Ѕ<h����ҩA�f����g��$� c;o�;�1��v�躥-Ey�e�p�%P=��5R9us�"�X~@d�g���`y�3	�pK�2MF�v\/ե��p��ό��^J4e�����%���f�i�ܡ┕ȱ�6cc�+G�:�Z��0x 廬�=ce�D8��a(���V�s���N��?���BZw$��%��,�y���\Y뮧�Є��Ԁ���ڔ�e��:�o���I��3 ��@���@��=j��7�{泻�� ��ͩ��N.6�H!�����c�<�64�B5��� a+!�MQH����d���o!E�=���v�q�C���f�y��D]rQ՘��QX�V=7��c�����&h���l�a�P���%��Pȶ���%��$q�u��UY���Ϳ�=���C+��+�p��Z=�bx�}3�����R���H�a>��r�~K8,4���[ ����~�6O�d5�)����j��ػΊ@��`R#$�#��东�y�Z��$����vӉS�l�P���G��{��Yx"#�9���n;�dQ
�k�<ԠI�~��:U��K�&~nٝ�e��<��&G�/H�y}�-Ʌ��f�V�C�\PGH��@�_�yr�M��E���C%�d�ni�-��A-��ďD�X�Yg�/��֠��#�@�;�>�t;����Z��=i>����I���-3�W�ePì��]~�s��s9m�e�G���Q�5�,^h�|��$U%y���r)u'��Ś�{�ҫ/cZ��8q�uk���	=H[Of�'RE��J%c�'Oeg���A���j2�w��*"�s3�F�h���H����'�st���[ix�v�H�v1�4����{	����$��:�;z�=��4��r�W�]O�椬ɓSP�Ԣ������V��Yy��Ξӿ�^SIi���K)Tmϼ������Q���Qgޑ&2q{g�v7��-��=%��S2�B+X�5~�Sɦ�P��ƛ�\'�M�u�~%�7v�eZ()�йl��6��@�o�W�O�N����r�ص��D��o�N�f&��G׼�qʯp�4�OB��Λa)�����$��&��>zLP3~������$���?{o�]�{�S���)�uR`���f��},�]�*l\��x���L`���z*��h�M�@�j-�bM�3��*{ʵ-!��P�(E��^���uem�����&�,`�cZ��P�g4C{���^�HY#�re�#f��x�f#j����n���}��[�����.r>��rE�DE�K��v7�F��@x~\}�u �)�����ڱ�n��?��<^�	>��qE�S��sd3�����إ=R-vPS�rekoj}�G�r���ĺ�Ԇ�dKs�k�`�MY3�B����s��.��\g[���!{t��1.�"ī�d���X����n`/�\��l��5������� -�A������ۏ?{[�j|� ����B�'�b�f�W�Cѐ���y�37
�Τ��N��Yzk�¤;'�zh)�FJB��������o[ci�Z&���b�"�L����^��,��U0m�S~�O\[���`���~�!Z�F�%6�AV��c� �"����>p��1G�_v�i�B=�/yq	Vے��u#=9�;���]�7��]y����{�͟��Ym+EI��a~�trܱ:P��Y��}�]��"�G�H
.�gƙ$h��= �_@�����'�$����b{�Z�K�k;�oŹ�j����&��j}�D��v�#@���ya�[�Qn�e�)��(o�.)�sկ���	G��ǆғ��1D7�|��;tq=B�j���r���!r�P�m�F��K�6��zZRx9"}z�e�YB|uk�R:�kĄ�2P��v,�Ц��aqm||�`"�����0!���V��ky҉�=/�Դ��!��i�h��r��Ɨ2�#Z�U���JĄ���Y���A�5$�H�܊�uG���tNV�ҫ���
sAV�,#wa�*���Z%�o�]�����1I�Y����Qt��xGy�v���U�M��P�	R��ʕ���<V��7�$xW�>���;�%�,�-��-]Ǣ��9|bM-�|�]7��bQ�M� �b0��
f���n*�G��d���a��a؆s��K�'��g^�I0��_󋓕�[ث���͸I���C���N��ma����&�� B��;���^^a�ZP2?�bD�V�8��38�;r.�=�U����Y�`R��~
�EE�
�#����U�g7����s�Qn��%X._l�eG�j�m��2c�?6Uʌ��cǩ8����3ݼ7 b��ϝ���P%O�[\gӒ�U<l���%��C���j�ZϠ��=��A`�0�x��Ԏ�F�BI��ͳ�/[��G����6zCkN���"����=��W��v���{@�#��+���GcA��#��X��_�{?�[L�AM*��I����y�(>�!+�SC'�N[=g�㈙�W�ͩ��j�����j@b4�B's��$�iSH>}��'���m�iI x0�~8·��k?�Ʌ� r�3�N�B����K��&�Rf�uowQE���?�$cl)4
�|P���8�]\�L�X����4���c���q����p�9Y�/�%0�����W`]$�?�=eSV8��:����r�a�v]5L�Lw���Wz��LP�
�dI��ǏsJӑ;����~�p���η��N*�=�5����=�V��T�rg:rp#�a�XD1�U��/�n}s�N��8Bq�]l��Փ?PʩK�\���۵ ��@][�8��f�5��H�� &�FHyѦX�ܝD�e�Ѵ�d7��V��q��՚PTX�*(�F�wg���vs��,Z�Z�u{Ӣ=mP����O�7ZU!�˾�w7��z#ܱb0�g��qYй�A��Yؑ����	$��L�� v0�k֎ 4��;� ��xͫ�׈���h�?F���ޣɃ�L_KƉ�Ki�Qү%92��h���}AO�f^��8xY�1ku3xm_e_���*0l��א� _��������(.*�l�1�0$fա5c��?`�
X�����M��6&�e}�F�3��1��>�.q�f��JH��9�HZn�����Uʞt�q�Z�\���K���/�|^-����*F��wa�Y�"4�y�\Glte|-�@�wQ��!J��v��ë��"�6��
-�)��
�T�J��X6h�]K;.iq�T�;]jſ��7f����'q݀��p%��V������ȸ䋗Q�Co;����|����I�0�����g�z峳�����k��x�0�:�����:�m?��kczH#U���[�04��L��c4��fFn��V��&l�l1��j���
�Y)Tw�`Kߡ��m�����O�
�([O�3�R= m[�Wƾ?�?��6�s�B����G#��n9�
V#e.{�(����i�/���p*������í>�֨����v�����EzB8�tl�+������
6	�U�y8�6��;���%�I[���ҿ� �2Ѭ�s����TBc�z��ސ��r��-��q�cQ�v���';=��樫����/����AWbp�q�&?j�vZ�C��>��\���pz�PD�@�n��ʥhi)�ܳ�\a(n�b�"4nV�M5����|��`�|�V��  ��4�wY� b|b��f���Ð�w�:s"#�A+�w#�@hא)CDE`���i�
��3��y�»�'&���M=~�@�<0hxk=�q����m����i��e��q�,�G��i	aV�H��&(�t^��T 2X�lx])���Qp]]�
j��&��=�;�}�����q[bI �>Djs{ĞJ��djjZ�fn.["kn�c�$�q�!���}��aX���J#�:\7&�b��CjW����QcNL0S���U[�"��@�[���~�B�(���U�[�^,��j�֨�s�Q|.��#c��m��:3� ��%��0g��Kw�J�1�h�����S��Wm;Y�E��'��J�n~4�r����e�V�u���ϽF@�_rPe�T�� d&� DJ� ��*H$�Z��A7�_U��7C��l&{�A(epև�Ά�b�S�̺�N�U�6��Z"Em�y:�eۼ�����\)��_�Ò.bd�T����lPXx�w�r7ݭ>��Ly�q�V���ܙc�c��J$nئm�(�+�n�����"ݕ��n�+K����ZD�5�{�ͷ�@S��6|��θ�TBV�`���BÝ)H��<��-�=���d6�F��МA��z���,l��34`%�w�Ymk�m~����Ƶ��F����� ���}#)��aj.���bxi�1
�o�י0��d5 ��)��E7�-���0@<ƬC��>�h��G�� 93�[c}|�B�`�4u?��b��J��1kI��Y>x�m�bL�v\{���XfpP�J�8�����w��=v~�l@��.��d(+h-Kx���ȯ������i��w��knLNS�z�:�z{}Q���5vk͓�ې�����=��ls�4�8_G¨���naYj:R�����/��vK���Ɔƈ:7�ۤ�hT��m=_���1+H�z��"��VQ�O�/�>R��^ain^D�NX?)Z�O�;��߷�߈J�	��3��4Eڳ���gK+
)5�T��O��8f�Vo"h��҂X��K��]��V�5x%\t�ߦ�&��q�]΃'W#+�{�W ��e>�R��2�1h�ַR� 9zw�jr��stz#�_��MT���L� ��	�)�N��B3���v*	߰�����y)h�B���g"�r�H����ʠ�/_5�#*ᩰ�JPJ;�8Q��	�Xv{���D<�ζ��^�U.<yj5m,կ����3�ꃍ���،�="UWؘ>��U�5k���*0��z@���_ӌA$2���QV��~7�����\!�wi�^�O�U�bv��
� �o��h���~!ذ�6"c �b!G�=��I��LE{	%N��ԕN��H��`m3��*�4s
GJ	��<�x�ԧ�J���h4�ZSH1Ş�Q=bsR%Q��ؗ���ԝ���sƾ�.�9O���
b`P�{C]K�)��Y&j�ڛ~���Rp[e�kJ;��j�(�C[Dt��@jAx,��[���_����A7�-a���Ĝ����|����D���LK�є�Na���կ�6�Λ��ĳ��U8"��iۼ
�esM"2���OJ������ �-f]���@L���6�|�����S�xz�'Jn�2�����s���4��Qr:�ljh��[J�:�f��ԉ�W���f"�,�SMn�\��"��Ģ(��;l��9h5��hy`�mLHZ�X�D�;r:�1�-8Z�=�� W!��Q|�R���BXR�ӂ�ܷ�������ݗ�eE��p�cY�{�{���p�1�;�
0u�n+beq���`���U�v��W�E���5�q��5e�^�y�����j>[L�#W��]�z����'yC�D,[8榌�1�)Y��>�6"�@[�t!ؽ��5rq������A�ī�ʟIu���0�Fq|�5DVkk^Prg�䞻;���*t���ZF���o'Ք���	�mUֶ*ʺ�!l���T4��5?�52a�.��@!�1u{ cl��J���0"*�jb�F@���~g�0Sy|Y��K;���r���%��d��nn=�OG�FUk�3���������.Ey�v�n�-k��L��M~�T�\y /B�5��VUr��P�w�ℭ�|y��G��l� C�`�|{��VEd!cZk*h��4��ul�Iܓ]_��aco.�rDbz�(X�0Q�cj~fR/v�|��k�d�h��9�Qo�ACK���MCEDY6��pY5全��Z0OV��F���t.q�'�,�X�%}��z@C
��o�}0~��������2����߬���v�/�Ⱦ��h1W�x1Hr�t��-��ss����{� �u�=i���s��?���n%��.ʅ�@%������9♅��$M�%/"Tv	.{�ƞ䤊?�ϻ�Ż�D	 i�F��*���b��u�[U��!��,�g�L;n-����#�r��jo������>�d|��~L���0<&Y�='}g�ʌ����2����J$�-�B� ����#i5<�7|����l���-
 ��a��L$���9����뷺���6��^��	���N>�ji���L ����`��G�ۯ���$`;�	�Q�KZ��>�4�\�~Az,dl�FR����HX����U������Tv�����e1��c&5飠fOMx����??b_�(J���0ׅ�:��UA�zo�(��Ę�?E�K�:q�N;7�ۘ�B���L$�:nm�id�����\�EXt���"DKbP�,�m��*Vܜ�Kq�O\�=���� �­�m�S!���|qS��b�^���ޫ���I���4p���և�8��Pc�p}��y��'�|��w}�X���i� y��JTb�r콣#�u��u���
�0t�Qj�fr�
E��<���M&Bȉ0db�W��9
S���ڄB�i��67@x����S�tM�u.Ԣ3�%s�3�� �Z]|����kP^�и(����T4<X�l�Ȧ�$4���򱎿��H_��@>{�D�B�fJ�7y�j�P(}+�o_�\��q��'�=�zÔ�%~�TF���û����^7��5C_�-aÏ`{���_GY�͊t4d�Ƴ|v1��Η��~s9�B �.�v�o$w��.+�Z)�0��K���'�0��?G��$��N��������7j(�?Z6��hS�W�c�Ty}R����}��+V��$���SAmDT!��|%��}�����/�*򵵢9p�sC��	&��̏_�A�V��?�G���2$Ʌ��Y�	Gw5t�4��K[K�kmc�*
�\֙��Y)P�F�b?��g�h���x���V�"  sM�z'Sвv��L�GA��Gq��w�	��G��!�%��guz��Aɚ�F�|s�4��~����_���L�q�Y޾������א|!��#�r��}j�`Z��K��Q��l��1ꉶ�7�ڡ�����v6�{0��u�5/-|q�fI�&�e�{8G��[a���XF�F�:�� ��ܡ8����_��^�����L��j¥��`x�0�ݖ�Q��0�w�ڸ�~3�:�5
d�����b��_����h��ǎ��5�v��6�z��T�2h�_FB�9���X�Ȇ�e���v�<�q� #�ؖ�����@ˢ�X�DC��3�CF>U8�]����I��Q�=Xץ "����PM^"�i��2��������<ƣa
� �^�s���k�~��s������:݈���\\�B�����������}`D���\)e*g~-xy�e��9O����L#i�n���yt�p�<�I�D�1�$�T���C�����bM�0��r�j�Xy:C�/}���9�:�C���݋9�!�	起<A���kL����>��׷mǐ��/����B�>*a��)�ͱ�ͥb)B��ګ��������f_�gf�8*җW(����(�䰳��R�v<�(�&t��
4t:������=鉝�[xOz�������֓��Gf�P��a���Jv���V������	?9�T���i@���܅��\b�[��T�)�'hi5�NK�wY���ƎBi.�P# $�L���/��	9����hRr(�f�a��@��&e	��XN��7�?���nl�gО�C��qcP�0��?&Ū´��K��TiΕ�1I��_�\������t��uD2�4q5���B�.�g9)�Hf42)1��Y�����N�' CE=�:n�&`e9'a~��U���/����ϭ<" ?�;z�v��=+�5b�iV�{c�B4�0�7qCkh\kUUs�-7������(�@ŇU�����Y�P���-y��me+O��[��ȴ�1>��C��\;�r/=N7N�̕���������́!!��I	�I�ǁp���H��<����b����L�?)P�tS��}Z����];�x��] :�s���H�OA�h����2v����o��O����F��! @�'�70*\�*�õ���3�M�l�^��6]��p#V9	�V��s��o������ ��TA�&�[Ix��Sx�
*�np�-��x�P]*�v�F>�%��:F	�9��V�w[;��0�����Q
'�?���-mġ���T�l>t�� �;)�6,���޴(��Yw����ӷ� ��JvX��_��9$԰�[	�8�8K-U��c
l�er�����������bh=V��]T�|�D[ܳY�[��D�>�j[շr���c��߶|cF
�b��W�D�Bbd:T~9<�Xјl�e����يf��Xd�	~�T�1O�sP�uA�������-#dB��R3�8�)��r`1|$�� ����pII\�4F�OӀl�ϴm�-{���a��7 �IH`�;j>&E�M�橎���������8V��d�{l0�FL���	�y1�(��Q�Wd�P�v�dPl��O.$<�5@�/�"��c��41H�������~���7�C��_�8m�ts1of���I���y�ߔ΢S�Ch��i����s2�U� ����m�U���M���C�/V��ꃮ�+."C�t�I�7y���w��8�� C{M��t|����a��<����ɥG��IbD�&\8E���p���/P��T֪�N�������_7鋒�t�Wq�Bw1��o�T.
�T� �mUp�P9�|���I�	W��'ކ�ӯ�O�`<QP=_O�	�y"��Q�Z��glsa�Qr�u�|�L� �q��|1m�aB�f����������:}lWr�!����Z# !��;0o�˯C� Q�i�]���`�H��6�,���Z�?m�>��a���<DsaA9(h��C�h(E�p&?OEI˹�������[0`�a|�O u+�n+5���0\�+�a��0Wn�4��@�o�H5�������W�J���>2:.!��{�m�V��$��{�h.�iU�%;�����f��?��]�5�i��L�z{�&_��<E+�6,V뤍2�k��Af.iY\CcF4^���:�_獿tR�}=d^R��c�`�m�~�\k)96~�lQQ�ug�����hd7�^,���QP��V��е�0z�s"\��%�2Æ��E���nj�	ݹ~U�í��ŝʰ�Z�\ZS�}����{xp���h��g������C��&q��@��Trc6�<e:eڝ#1�:R4�!�9%��S͸O�'���8�s�j�c|��2�U6r_�`��~',�5*\}דm`�D��X���(��c˧�:��x�F����T�����!��:�e�5e�Lq�ꨤ;�̺�i�/'�3ѭ�)��H��u�h�j�G_-%=�-w��UuL��8��}5�r|��F�Z?�S'�A�^�˧���ǖZ�!9��W@>�� ��A�8rnu@�䌮b�������(�֜Cw@�/Q�f
'#�vҖ�nB(�@B�C�/�vR{
������Z�
�IF�k-�A�E�Υ�5�9��x.w(��L�����bT�E�k���,���p�H
���Qj�C��nʩ���&F�e�8��:
�}ք2bˁ���7�����tY9�����ُKQ���p*� �=@!�氟8��A�x�E�]�w>8�袋�1GE��kܐ�5��d,� K�.�n��5v�ds�pz9ê4�E�56�-;��;?�[���e�)R�I�c�9��g��o�:�<�h�0�n�8�K�Y:A����/�gƩb�qnG)��4"�o� �Ӳ&r]��}m�0#8\`��W7a"���Z)N�0�JG������S*�%Z>t��Wg�A��ivժ�O]O��� oթ-Cw�9N�ȡ�۫G���@PbD�ԗ�\JO5����7��`b!N��/ZM$�c��x;�߹`T75���U���LTA���\�t�b��%�7n��w#D,�!��,�1�am�v���� j�;fL��QC˚���a ׯ�@���: ��A��;$Dɡ&q�xxD!���~�N�&N�	�D�/l,$��� "`�0`�(~ϸp���W��=u~�+#�߭��I�`�D�ˇ*��{��^���$ی�L�m�,.|�4L�rk�U|a�G�~�������z�=�D�W��є�,Ng3�}����>�@}^	�t�
y�>4鴘��W�>,w�������މ����"��O?�� ��Z��t�u��]p�scK*q��f�2)ǉ��B�ׯ�t�H��fe���3dT�7-l����Yr��ת��ջ�� w��+F��ʡB��n0Љsa z9�n�|����eg��3	9��@����;��^���O�������8�Q�������W�����fϔ`j�������g�������H(Ř&d.������Y%Ƌ#��)��e1�f���uҫ_bO�IN�	n|k���K]i�<�B6�܋إ���UhZ[��g����,*œ�P��D����+�x��m���|��pI:��X��� ԠWV����	��m(]4�۔6KB��(y����mC�<v���P]��o/:�h>�[bK�� ��c�G?�nPu�/�����8�;���Z��FW=aBצG���xBo��+�=n�qEz�G�H`�[Jd�R_�w�-`ء�*v��<l8����d����E�u�H<����m�OhR>�4TF�)�@񒗪C6�?�W^t|� ������=����F���qr�m���D�Ԁf�#,�"rڽ�(ۈ��Y�A5���V�8�,�o�-dY�jC������Ζ[޹��ac2����<��vy�ʰ;shIq���Oh�it���f��v4jކ2`�2u�cʾ�\����6:�H�������KQ<C�t�65JO�t������wXz֗�B��,�=3W�>�1�Ձq��@u����)������96�Gա<ս�
]룰46s��}�_2�]o��G�u����ܧ��`�#OR��*) ��ld-��>�/ݛ4�����ge0�'*^^Тi9A�^2��?5X`�U��J�]��>m���d���[�4D��Ʋ���#͠����K�no#6^3����E�/c�F5K�)KW`贷~A޿�/�mʙ�7��U��u��2��0h�xs�+j��]�/�����B~�$u��'�WE�".� �3�'��r*U�م"̟+Gz�GY��/�-<YKY���^,�e�,n�R
���)Gj�G�©��v`�N��s�� ��Q��>��6��(��АY+I3�T�f��r�x���Hy��SH�75�z)� ��ï�-C�M�bE�3>i���¹�X�	����`<::�m&O��XX�LX79�9K�����G��F�A���y����-k/)㎍�l��
�}L�O�e�o<Y˷�($���+���h�I;ɫM��Gc�r4�ЀO�{����>�[�2�и�mI8܎�3&�3x�ʦ�tX�ۊ]��"�D�r
�Ud,��}�~�vEr* �С�Z��X��oy���i"������+�
uئ���B�3zK��1�l?��m���3�T�ԭW��kJ̪�'FT�8�J������������_i=+����2Qq#�~��zP��+��Ne}��lN�#��6߶Ev}�8C&�	mV�Q�T��RRwJ�s�+Z-�TuEy�_�d�/��clE��;"h9gf	�f_'���)�D�E��v�k����UB�~6�~&ȝU<n�t*�(�'Q��(;s�%A%^VW����l5��j��84�<�3c߉�D;����ݳ�6T��cl&�4tB���7(Y�d+d,���&��y�h�R��6w�f �ސx�@���)L�x�R$����txE4s�}7�T*eW����/�]�����E���.�P2�L�$\W����g�I�0(���ү<n��2�ϻ�Y��3<��@�EN��������᧱�ϧj�ps/X���:��~��y$ȣp������o������ԅ*ٚ��r�Z9wyޤM���7;r,����4��<)�~�~��=DT���=��/�"�ː�"�u��N�� V�bI�}�X��Z� ��I�"�6�mx�.W@���gnD^{ �Z��M���8����l*նRsE���鎚o��m��&� �tҨ�ΈY���#$#o3gu�����+͵6��	��� c��=53�&	��ō�jf��!奔�+���zq��` $� ���Bz�>'­E����@zkH�'ܓ<t_T�;�~�c�	?�Ct��A�UU;����\�8̩9W�%�w�''r��i_PX&kn:���ӞB�qm�}�9VK���~s¢��T(Ī�>�_��w�]�l_d�<Y�M�,�{�ng9�R�i�s� �L���b�qo�����跶Eu��n
����O#��f�yJ��_).ϙ6�+|�O(�1�ͼ�Pw��lO��/D����$�Ub"X�z��tO��1hX��
��g�6�S�e1��
�u^��Np�ĥ_�����p�n�.ό����J��4_�zSExf� xƷ�Qd72��ٝ6h��˼ �9o<��\x�X���4��v;�zоK������K>����X�܈����s�����E�#�)�ЎbJ�?AZ1a�߃��K�B�� �LOc3�� k��?{/@{O~ ���`5��P�ԓ���Y%�M���#��Ɲ�<i[$�_Y�4��N�q��%���;�/��o���N�RFEm��t�v�Z�p��A�8��{���)2��h3`�gp��+��9�fլ_v�z�ur��	< ��ɭ��uL9B��v΄��F��Ʊ���_�?�i��g�L:�Y@�����3^*9�l瓪����eX�G�,��]�h���bt:o�d.`>�-�	t{RI�o2Z���Uㄪi���Hx���/����y�=��	�MV�>L#��ԑ(����z��j��}�
� A!��s� hS���p|V�16�����P~
�򅔈�~7�)����VG�.Zl^!G� )�ߠ��6j�]ە�4C9��2�f������B�c��s� |�L�]��˃B�y&~��L�B���`�<���s�^JT~�=��H]�f���'�)��j���H�\@b]�q��a��<�SB=��K�1����{>��=%pf����3	���DC��2�EA+ׁ�z☝�8n V��`�f��H�
��7d�����2�.Н"�$�Y�T��eN�^eapWJ��p�i�j6%)�,0²���9\՝6�-%�(g@)ҷ��R�\�lD[��4ΙI���A�Vw*��-��l�Z4I$�&9��D��ԥD��gf�O��b���k�4����瑙��Ih����5#vi�ڻk'�T:��X��{���O[�M���<g^�5
행�⺤y�e��y&`i\��V�뮚�9}�b �+�0nҰ�MK����9+Y�U��/��[��.}E���M>pbیI-dyN���k��s�x��!zd�D��������X�$oW�n�}f����y��]�
�l\�����2G���Z�p���(x�K��|<��V����}�\�x���l 9Q��#;��^�I�V���{�,��eK1���md���� ԩ��p}`�n�4r@���������@�A'U�[Gx����5
��co�E�n6b ��>?�0��o=X]}�4�3<�l�(��4����!5h ���9���$S�Z�H�¦�={�Ri��rΓ�[�"����w����T��M��*�'�|0��^����Y��5�_͔�&c�����Hb�P�0(��t��ͧp�	��;HS �/�J��'7�?f�N���<�7oR�-9��	I�fk.�Yq �����mr&�� ��%إ2�����2r#�~��@�ū`b�iV|��o�rַ;���8C$����j��e�G��JƟ�Z�0H����?��y�멦��h�?�W��&�Q�JmZ]����>��$4%�q��|@m��&�aO4&�4 %�r�n�Y��I���b��l�Ơ��񄂌��K�м�'��;~7��ơ��z�ɫz���5�U�,M,���<^:�d�fܴ�a*>�*SXE,�-y�O���u�zz����A�=9��V��5&���E�k�A�x�������?�H���yw{�@_�� ��x3�A]�ٿ~�5D񖙬�9�|�O�Hz�|g>����|����;��Z���bJFX���a�As�Tm��~���c�p�9��i|®�}�����B��S����eN�"������ؘ�Jj���|:-0���$�V�P�=EjYa�iy�?	~��o�r��ٟC`R\g����f���i	���)�=�B�'n|�@rz�r~ο��F�m����eM'�S	����c�(����!b�����gK2���n���;H3�s��>�-+L���Ox������n���~��	.����@�8�٦�!���A�X�B�ɌC���]kqy�Sa�]�Үq	8/9�?}�a`�=zՒ��}S�3�����������|��|�=H����|�p�l���rH��R/���:�/;Ӄ\VL�ߐ*��P��x'�R��5U�34Ax]ϭ�P�?8���Tb?�!^k�*���d�9_Y��4�.�� D���% ��#��f��9Xdw�\8-C-�ϵR/w����0陿���|���f{���8]��~02�'��R{�2��V�R��7��k�R4	�3�#�	h�8ÅH��`V��?���U�{67��2Y
AsZ��II���\��ϴ�j�_ ��������|^��>�6 ��K�9���x������l�y��7Ӥ)]X<\����	+3�èg�űX�m<
���R�WLV@��h-�ad��JEM)}s~��O�tĕ�J�.�Rũq��N\��À�Y���.���hs�w�Z�b�@���3-:2ޛEF^�^wI;��QB�9�F�`y%ց{�&�� ; ����̤~m)!^�0v��>��r�<���e�G�h
���M5��w�˶�1Xt5�����Cn>cf>!�+�����ָ��|5=ϛ��N��M/�s�K���"�����K뾝�;�'9��|�>����t�p�җwu1�������$�G�2i�A{�_+��a<�V���b7����~��Ir8�R��G�j���4=�v�}�$|�٫�)�H�����e�5r���h�t�$s�A˙�2&ֿ6^(d�m8v~��T�V4�6���#�[8��L���DF�yQ�k��l{�!/����ٴ��.�p6�b�t+�����)�p��ax���T%b(�Q;��i��s֪W\��+� w�h#NZ���4?���E���d&�M�(�XJ?�K迫�ё'T�s�����2��"m[�����*׷,�����=]h��*r%	J�D��f�&�fT��h�����$@5��2��O��6I�u��/�+�>?�ڏGN$�w���]�K�./7����rg�V��f�m�8o�J�PN���� �x�^�Ԡ��o�Q��{�����f��%�آ0u��` �1��ݶ!Oa\��Cp�jy0Τ��n%�t+�\_�d#.�u�Y۠ʋՕ ���%Y9�&7�����or�&ƌ�I\�?�L��8�����%�>���˒���ώ�m��3)��0n8~M?Wwi�X?fl	o�d�̡����l�껏�k����{Y/�����z�?!��9�8�E����C�4,6�d�o>2�n� aMށ�O���ǓS3镩�[�{iN˷g$PY�=Q�����M@���A]��+A_`ԁ1�J���
A�����H�PM�4�Q d5�#�m�q���L�(U�:/?%W�Zp���5v�*��C�P�Կ[>�)�˶�L|�q:�=I��6�T�0�dh{�/�[��~}ϙ9����߶�U�B$EB|���3~M��]�o�ڟ�l���:�{b2�ޥ1���ӝm{�J���d�/���K�p�;/��:� j��,�~w���hN{�bi�-����m�,Z��G�\Çȁ�P����IbD�"1F�R+2����wf�QKk�?���},7ic�f�ۃ�Q*��y97��Є��-W&h̍�?����-�/m�~��ê�U��%�档��)؍g��v�8[~2��eUW�e���w�W<��N'U���ŮI��P�4��I�����a~s�Af:u*��IQ�����������!VnQ�A�4z�4��I�-�Ap���J><q~w�(�|�Ha@r��2����ܢ2�����F[�R�ȀW_��d'��$hȗ)��&�M��� Qް�'��q��O~�t��R$�l�\D�:�BMY_J��^�]^K�tI��P���Ǔ�>��0��6�+le
��Ok%�u�>�l�vQy0G����i����V��Ko��u`�!�ަ�&�m���dcfAuE\-Y�nͿ�.��J�k0o�����������d��z�����.b�H����0{����.�y�b?����%�[��"Ʌ�.v�ۙ/����n��G������Q�A��y8�"XD��U�;��"K�*�����,I0�����ۚ�y�a�`�A/\$p��#~��鈲lP����08Iv�KT�
���#����ef�&�uk/�xh@��k��O�՘�S�~���q���6�'�h&fu�[����є:x`�!�Jj󰷛�54�aE������G��/���D
4�^��O��a���C�����N�p�f�؊F�
0A�G6m�]���4C��K���$�3屺G����G�zq3=�X�6��	���mR+�VV�#��������^�&I��R~y��I�%������A'��y�-�!�Y��쩧�&jЇ�"E~U,�}�����Uj>��m��$��ӰX�O�Ӡ�s�,�DA����7�]Tj�k�߻r7"�����b��6O��,+v�v����Ŋjm-�dmeY��ƿ���[��$>��gX�}g�M�u�PL�t��L����f�0	���lz%�ޤ8F汈 @�c�}=⸒���W�C�����V���D�����y���T�2�`y�[�_&ٍi�i��L���tjfy��v% 2t��|�\�����L|��ҥ$\��UTD�{�A��J�N+�2�{Xͤ+�]���W��ü�e�eo\v� :>�_��0�%���@(�-��VW��٧�㊏��!�w�݈w�#�Ё\e�# �y��,���&�b y�*���6�ፙ�]9��N]���r��E��]�u�_� �����L��?*?Kb�*B���������kռV~���x�}f��g�d�ƗYm�J~��so$�pqU򷛪��T*��~�zkFj�\R���eo���ű1�����?�,��A,�f���@HF�+��ip��PE$"{�#ȼ4��K��g7�]���Ŀ^	���m�L�e ?L�z����YJ�T.;����{`{���#�t9��V�(�6��`��d�0��`B��*������vs��=��et���_�z?����W��E�rH��op���glXO�>�P�0��X_%$�e/C�"N��Zױ�ѱ�el����.,�XY|����S�s�>�)�շ[�W+���Csʄ��>Te���'��|�jYoVX��U��F�!&_c)�|]�Z�w�H�k<]{�X���?u�W!Q<��Wy�?�ʋ�[�����䡕�xM6���'���^�쁑v�H,���u�����$��4��0dΏt{�\��߯@�o����2�l&[��H*��H��N�Z�`W����u�mf9y�L�qZ4�C4��FO�r�/�9�E�$�z���c�k��G�W��`�^g�H��m��)"�4��v1�;p�l�N@��(
cN�g�_ם��f�;����^f��7,�=��	Wr��٣೭N����,[O|Rѡ�w �(����@��()�����K�WuJ6Q�;գ��S�� �=�NH[@���E��-��_X�]ұdg�mx��1yZ�7Yb;����P��$=�o�:���a�"��>x9�	Hg��g�ǘ���
.�8I��A�"r)}oa�C�T��h&��Uq������l���̥ȍ�;7����Do=!{�)�T5� �':<H���]�f�:�.�Hz�XG��YJ�ν����(8f��o�A$:m1�:�&��
�y���Z{�R	VmEt���P~<Z;����#�%ӎQ��Ŕ��f�Ȏ��h�?��ێW�� �N�VAa䝸m��5�\
Y���:�,P�WRa� �,P9j@��[9x�`�����.�v���i�����dc'Q�U/Y/�gj�r~�風�IcA���蘗��ɬ���Z���9�[��1�'��'��A��)47�g�����Sx��DI�AN�唘ÕqmmTv���_S�QC��芦Fw��ቷ}%�lDǆ�𨊾�T��N����xX�@,�c��b�9�Ǎ&^�{y/&�'�D�p���?��ꉺ��Nr=G;	/��d���}m����֭n#0$���f�}<���3������*mg�ȅ-�:��e�:4�AT�Yk��`��l�5���A�)�F�傞S'1�<9r��1�.{�SE�ğ�N��DFE5�di�0j�[V錧�#�+;f�T.8&ȍ\)R�C��3��D,\7:�?�`�Ş�Q���W����� 6~ִVϺuR*_^�E;fs�� �)�T',��PsU ]����2w-��y!�.ꍓ���x�����	���mD�ўeJ��y��H����I�ѥ��w���I���������-��~��D����2V{����Vw�6O�ah:�ً���)wR5�P> x�nM<�4�ܥ�6<��`�>�n��0��,��ֻ�Ӱٲ�cf���X�K�	�!zʢ��3��ʴ��Eu2��:VR�f(�C��6;�y:>=q���3�>�:�S�^�z��*�,z�LW��="uM����V���z�zH��i'�`>q?��{A#`�W��e�4:�
���w���Y���ߒ�I��L`o*u�#ĺW�'L{;iY=0�u$晨4�a�!\t��J3�?�W�ҭ�����Vm)$Hc�V�xA��t�rҒui�ͿP��A�7��TL�0w>ex���؛�Mw,g���7YLB\z5?<��R�H�e"�X�O+6ޗ'x�^(��"Gnqg��\���rS�l�O����G!`b�"�!�(ˤ�^�޾�^L<�nl���,���2۾�~�x�}N�5������e��5��/,�\�.V������Fl���w΋�Z�����p\�������%���R��yˍ=���a��}es��M���
��Ժ�|Oo~:H�i3M3�FW��Xmɍh�d7YK��{��o �ߥ���9�D3#��wS`"�P0]�HpI��.` ��&�Q|��Q�AR�`Q@����iB�i�3���OYG��y��!���8j���h�3�P��PA&+�L�>�L�wi�[��F��_�)�L�o���7Q�I�[���i멫��=�q���`)p^�����"= ��m:�=&��a�)%&sT/�I[
���f\9;:>�~��-����^�(����������xtJ��z-
����p������u��y/�B�O����Ѹ��ʫc y�W�c��������0ً�Z]�sNaҼ�.{��-ZS]�-f�6,��t��t�<*�,=��[犢T�����B�'ݪ5A�4=*��16^��Q����t��6�,��E�S��)Nβ�mp�u�W��Pz�?��ݡ|L���/̅��[aޠͼi�(��>sg��c��;�Ё�����-j��<��,����{]~75���$�A<���:��!&x�V[bRƞ?�T�)�}�!��I��&s��dr�;�̞N�9%r����+#:�� ?���1,)~�-�Ho�+�Y�'�bv��7^$�UfF3�Z�Ҁ鮙m�u��юF�J�@?��V�\z���&c��O	���U��z.����p�*_'��� ��5����ौ�J�䗂����y��F�۫�>�������H����əgЇ�m95�G�u|A����	TFwz�"�n!���4a`@	O|G]�SX��,�-�M��l���Br]lcr�j��]s���]������S��7�}�
��B��y�?�4�ϔ{}�L������gL"!� Mـ��Y0 ���K}F��,)���Ǭ����{���~(�it�������/LtD�*^'V�˄R�s�K��yEc�e=j�������7h�xD{;�<ۜk�n�%��>q�3pTl����`@���N��	V��,�A��R�M�,H(B�M�B�ǔ|��u��� ��H���AG��k�=y��3=���7o�p��X�"իݰAZ��^F�y9�9=��b�c>[69��SՉH��Ҡ?|�7T%`��'�s&�˺~1�D�vV�����8���N8�32�m�L��R���A�]�O�98h��(lxf}H�	�.�7��� �W��}��n�Y�<˘�$40��Y���i�"����I@��~)F����q҂>����#���7F��,�78�ضq����H���!���V�~u�o�O�C���@�4�[�]bY���"�8PAZv:ap�݀x�<kA�mTt�&,fU��l���U0g��J�=@mru���˅��#�����/-�إc&�<B�dh�|E6��V���g����2L<U}�B����m��\0Վ��nK,�t��.��γ���&r �u�/c<�st�_r�4�)���6-��<�&(Ni1��^B��s�mep��}��2jQ�]*��!72,ɜ�-:0r3���Xn?OS]ŧ�i��ˁ�����������l��:ӻ2!U�Q�zi3T	���|=ld�ҋ�h���=X/$���X`��)Š��VGזw��q* �,�6� ���Y]
П_���P�S�S�d������Iu8X�`LZ�dл�MP��V�C+WC>#̑�`��x����B�9L浇J@L0p��L�*@ۤ��X�J��l �O�+��w�)�5�&�ǐ��g����,o�ё�}�<E$�W�w/;8�d�#�j#�(����W���r	����\���G���H̝�s�ׇ>~�r�z�7i����~��
�{�%�
4N�{Uh�47��������ʤ�\ӑ�uO��e�6/�"�Ȯ����	m��+�]�c��$qh��Mv�T�sMjV��ݣ)�Ri���G��<�Pa��4C�ꐠ��
wWΙ}*��'��O��@�F�b�U:�5F���γNta�����������WjX�t��D��#�X��NS��
����3Yo������PN�y��GN��J&+���v���fa����^%/	��^��qi��m�����/�ψ���2A&�t+*��yT�(f?Ur��8y![�q\�g��e|�"݈;ю��FLs�����߆��6��lh]O
�FZ�/�|���Y���- 
���VLޢ���%�J��%7�X��nޤ c[��d����Y�CN�N��Ѵ�Ɍ��Ǘ���)����Ӎ�*��0�N9^�:�}�Gw�n�Sߣ7񔾋��l�ƹll�Zu��QI�ι:�/���:�l6ϫ����k���/#�I�̸�.�ˇC��X����.�
C'J]�[&�B�C90�燽T�vO��y}Ӱb �)B��I�J����n�<�ÏטlI���鑉2p���c���ɏ����r���^��q�G�J��+p"�olJ�B������RG�/����C�D�6+D`��﫣�6h�MW�n�۽�8�aY�GzS�A��#ϧ��v6�)J��yp\-s֬�4v����IҸR :����r@�A��Kh�@��b�2���7R�*Gw��ka�%�a\N��2��Ó5b�#�ќ�} %'���"ؚt-l` �n�I}�׳�A@�MWB_�3��@�փ2�lX-e��4������;'ʒb}��r�%���+�"�Pf��ݛ��u�3�&�P*'���50�n ��er˝Fw�+'EI�fg��k�eX���g?vu�e�6+�f��@�P���Z���WlJ�{z��61�l�o��u��-$6(�4]�\E�}�����Ծ���ெHlkR� :�Z�q�.�+�J���C:��d��I'�qt���d�K`���N�p�Rp�+"A��+b�5��Z����ʩ����
�U���1�Ъ����H�ȷƩ@C���_�s7܇�}nv<����1$?�){F�8�����>ѹf	çg����я<3l#�S>��y�75c�u�JҵpG2es_�c�+���l��Gǳ�4��|+�����*�u���@����`���K��f�O[џV`�6�T���4 ���!��<��_������)oU*�i�&½�|-ǎ�+�Xŵ-s��rx�:b{êM�����1���Iֶ3AX����@�Rk�����%�-x�"ڿ�j��b[��,Z�W�Ϻ��V�יF֠n�.ׁ%֍�A$�X�l�r�K�z� ᎝��Н������v����H��Հ$e�.�֯>r����O���H���R����]2o �:#��{] �N_O����BE�#��ޛ�(�j���S�&؎z}ـ�ˎ�5��('��bo���sRu�O��u��Rѧh5��s]mG��#��=�xz���H��tI�����/�D��$U����y� (}S�Z��4�9�&��M-^�DN�טt���r�"^�z' @+.
t?������R,��r]����]d�Qo����'-�&V�*9/��?K!06cH�^�d�qi�r�5���_��OKւ ��#���n�' ���U���gô�h'Á��Quۋ��\��)��@$=�����.�W�s���<K�{�\�I��������S����_9�-v9�y��`�3�����)GF2�����nV�x��jc���F���g��<�x�J�I�Z�uW�?f�_�I�Qo�}t�\����w��rhP�B)7�g��@����OmlhJ~�mB�=�B��JI%S�A���_���eA��M܅ˌM�����zG��+��.j����-P/��"��[���Eh7
�ܺ|��<�1-���o\u0p4�o�t|p x���D	�i}d�Ƈ����<���'-�HF��#}�D</������o���n�����B�`^�����ւ7@yPm�J�4/�;.�u�d��������(p�..
h��/hą?��b���_G���#�qz%<����z���l\Y�*9�xV�� kSh?����Y��F7��5��9����@��,�]VC��GbLl�����3 :���V�k�<w�k��?�<b��n��R��=��.
ݳ���n�n�4F�^ZB���;���fG����sW&��(���Vy�>�U3ź���=�����혊&�̌��ڏD�����=}bZm28$�z��*�C6.����]�����~_���ߕٚ��߉�e :k�:Y�&�W䀷��4j�� �0��JIZ���ۢEgmYf�FwR��m�����
�7�sԜ6�Ƒ!�@: ���KA�#�= 9�)��<>�`��Ϧ�Ҋ_��H���z��D���a�V��$>�>�|"�,iΕ���`n�q/�Em�g�]D��ۜ.���~�:��wm R��Mah���Z�1WBw�I�S��Y��u3�^�=��[��shkr��;�T�ݜ(�k�6��>�4p�3:W�����q2��/�?��D�8��2��������{�Rc�)�inI7i������~�E�x�>�O��A��n�P�z]��D�x(���Q��n��"R!�/�
0/x6�Y�����{�?G�'�N��A@9�����;�s��቞ )�e;R��D��Zw� ��0�s��
z���ס�re�PWL|�x>:L`��*��\�����L͊��a"��G**n��X�,�z`� c��P�4���2J=߫	�9٧�K{~���ջ�'�3���.8fT��&󠏅���X��>�u��/˶>8�nrǕv��8�:�a�>1�?�I�T�s(��y(f��;ء��ý#�{T�݋����)+���2yTb����V`$pӃ͜=iP�KOP��p�mz
}���w!6�<nvv��~��ْiPC|	=(8�$�V�9�`C��CP+�zJqjZ���,�����ڲ�1d�1Gj�p$��!�����R�����g�W��GR�v���f�;�����ț�/V��j�J]�xA� � 	�jˮA���y�s�NTpv���o1v��!V���@h�x��1���%��3Zrj��8���o?Z��18=��H��ՐW�7
K9LE`��(�a�l�o�<��4���h���h����]j#`��)*B���X d�e���R����K58`���T}�9������<o�6]q��O�F�_hgqUI��Q�=��L��߷Teʫ#_Ƣ��c�ڰ�x妒[
�0��k��r���A9"�"�&\w�t����t=�~��&D�����e5���M%eMl���G6�S�H�z�^�ǚ�^'8�Ƈ�#���G�%$�u]A�-�~�K%?�n�\O��2f�Ϫ��/̞�?��[XU����K���Gh�<B
"��6���ރkXmas�o��������.�y�
��rJ���*��[�l��]��lx%�UJi_�^���$I�.H���K���25��*�R|c����ܤ�9��C$�Ad�� ]ĎV����d�/]\ڵ.;���`/��Tgg������(Δ͛�,�L�c�F��ޒ��D!���}8�x�|���E55V��!m��዇�~���p)��17���[.ܪD�ˎ�4燒�`�A�#���~?R;��� Y������f���JL���d�S㕠1K������ԋL&����hy{��=BƦ����"�Q��:�����IWhDE?k��j�2#�Z���3+�?dzB�n��������cB���l�>+�9�^��gJ�+ �	�'sX����T���!N������J��h�(�Qk�-���̷1q�r�����u��<S�`�z�Ⓗ�-Ⱥ?Y��Y�;�}F�o�1x�$д�
yd�pҭ�u�T��چ�֠f��ߎO�E��vM=�pܜ r���>�S�A�R�+�%�Ayc&А�Q-	��$dG�/PM���R��d�Ih��MQ��A�^��Fea<^����;s®Ӈ]����l|F��W��}� s����"�Cw�sfX�����B�A����hh9�ڐN� ����"��9p�!|$fډF�����rIpA���&Y�ď柧�.�혀d�K:�)�n�2���н�1�4\�ܭ��A����I�J3 �YYCQ��A�͞vUU�����y�6�?����8�}�-"1ͪ~(�XOJ��Ya͉���(�����ڞg���,������9�l��a�2�
���d��;�?00�ou�n؄�)Ь0���,NO�k��I1n�
x��7���@$3�9�a�>���I7���Z x��^<�}W�FṌ���W�RGĥ)*48��5~2@�}���Xl8�����+�FG�>/�Pq�A��e���\�Rw���ַ��g凕3���v`���@�P�uġ�����Y7��ΤIP2�G�� <E��2=xĠ	��=�&wre�X���a�3��5��) .���O � P�G����?��y�����fq�����A��3�U,g;��gŝ{5'�:�����c�C�{ (�n��!�_���x91M�g@N�Tx����h�Bn�W�/�t��f����=���w~��Q�
��ch/w���Qs��C��Y2��L8�����=��i��!{\��>��B�ۂE���6������8>d�5���?��kМ��QsU!l���r%��n�~�;�Eo�^�G,��9{%���q�uj1N�|��ٚ��n8cBUw��(����H��XY3r0uS*���Mn.�ҹQ�=F;"e.m7���^�#���^� PĔ"�a>���{�e��ې.8���WF�{<=2��!L>xNǋ�W���m���^82�����c����
dRΗQ]!�ď6b�<u^|誔b�ɶ�ɩ�c`�~��$c*,ݑ�Z]]O4��b,��������{�p2���ph8��I	��~[c�r��'�\�&�w���*�kh�($t�HpȠ~AފI�E����������B�Ip�}���d/�����:��Rm��F�ŒM�����!/x���D�z3�������@���/�Ý�k0��j-�8�1�6��[�+⌸�Q	���3I���n��sL,�*U���jf3�0%	��K����\_��������K��!�>v�� 8�k�Wc"�٘|���6nWO���r���`���%��;uE��X	r����:�(���^���������Ç�iH_
r�$�ats_���>��]ۙ�=aw͸�ĸ��dV�u��߀��zWۅ%���.�'�l�x�eűղ�2�a8�x�Hb
�Њ��Nԥ�@\���{>��}�E��X�?}Lp���C�/��o�[jn���i64sK�I&��	S��O�G��Mʮ��ׅ4���.a_��o�8+C��忝���&I%BĦk����W�-�ƥ�RYTY�o��\�����,�[�]��E%�E����Z6�ik*O&*{�8��z�3P�.���5�-�)�Y�mٶ���˯Z����f��DB��!���r0�����~h���
Y�@{���Y�R(�T�}*�6��|T����� �J�Qh����Uѳ�b.#�'q�ƭ�-5@6E���Z]���j���%����(� H�7��La���,q	�0
����:Cߋ�,6�0�SF�_C8��蜺��D��N�7��)9@��(������+ܦu��sd����._�ͪ]v�����ۜ�n���
C��J����+�)Ӌ��p/a������ޟ����lp�����!V��͔��"�����p/�_��fЄ����v26�����͆� 1�5jXs�bN�S�� ���i[�c��Nh�Q�֭Wp�8%�*NN����)�Fܑ��И_sr��E'ng��|�q�C��?g�+_bt�1�4�|��n��9&�6�ؼش1o3����<`��ɤM��]T��o�b'���㹺<�2@��	�DX�	)�9Ky���Zy/�M��m�����|�JUłb���
�<{5��&cO�3��<�i��'r�45q�Et�ȸUc͕�X���D�$�����D�y�w��y�=���uT;��d�*ݾ;>2�K��y��+���;���@ov+������P��e�	�e�^Q��K��ac�r�4,��E�[N�סd	D���2x!_ �Wb�՝@�ֻ�����#ܗ(�
�H5:X�e'�����+�+WW���v�[����O��c�VL���mH��1�va�4y��$q �d��W
su|�h�A�	N��t�G\�[���`4���e" �K%�5ߥZ)��Mٮ��dʣpC���䕣��a��>��� ��L�t5�?�A @^_��4E�z�.��R���c��Dg���q���6�&��c�wa�ˇ�dץdiW��V���\�,��������&�%�{����vxV�Kp�*��� Eٙ�ߒ P�Q�c��V�t�$�ځ�CB�u~eU���B`��+z����\jU�r�����? *�&D�x)�Vέ�F�5,q6�H�1��t��g	!ֺ��o���NΫ�鍚?]��x�I]�{�B�+����t��U��MD����l�N�\j��g�D@&�O��mp�?|��|�.�؊h/Z	шp���F���s�����r���`���~�" |��#��u=���ͬ?�ywl��u�s}l�o聾�pAϥm����g�*&������f�f�e^��5M�s���a���p���@PM�l�SטWk��S!�f��L=a��|+#:JD��G����`c��I�h��<$���JМ=���nyʭ�x0ڴx�v��@��g���w©�	�\Qspq�AI������:�!��[qt�j2+��������7��GX��򿱷֩6���p��-߂��-᱙2��i�hK�D�|9T�ڵ���_��G������H�G�sv\B����H��."N��v��X��U�tH�E��)p�Nr�?[9P��`_�V���+Xq��i��zj��^�8�j�⼠�[b�.6됛��ǉ��nz,]�*{�������p�@�]Y������mh�y&�?����O]SQJ�k�o�t�|:�9JOj���F�[��L�V/;['��s�*C��)�"W�M�C
�i*�&�p�ztu�R�z1�˂!��N�T����S��o.�6P��)A�];@��=��V��
���Ηi��e|�����R��4-���,tZ���_6���%j�P����[|�㴌�mB�mvBC�%qҠ���4&\��
���[<�<��uE��E^�h��5��D檭�{��b<8�MO뙫i]�N�L�ʪX����_
 �+�4���k���`~SK !'�]�by����4���s�N��u�&5��v!>�����y*Ǧx��a���/Z�7�h�`�/X����9s'���o�ݝ]�b.��ڥ���Ϋh~;�����8����g�\�Y�>�e!C��?�_R7&�n4K���&���1�����4��D��4��S��D����S�1,�IJ&��d�Z_�D2��3��VG$ɼ��g�7B	\*��sG��'��$���e&.�Yi T�9ㅬ�B����� h��Q����%{�\a���![��y*ѝ�1 ==9a�RR��A�Ұo e4������M����9��hՑ��Y@���o��ù)���5'E|c��5��M5ؒ{��/7j�+ܲ�wi]}���W?*�]P�0]��7�п�� <�Te/�ͳ�N�v�Q,G�
:��_��i�fp�a���q)G�N]��n����k�w���zi9�M��������S�6�N̵��q����& ��&���S�G�$6�n�H������5#:�E���'c�=�ül5l����A��3<q���D��=V��1�[��?��-3��F
�?_[l�d	Cs�	.��H�bu�p��j^���D/��˰�����l�uJ`�"c*CKn"���K�.	��Eq��P�s�?����4fXQ�����n 
r1��B��/�9�� �|۷n�ܸ�?��5�n0:�r^��v� ��9]XD j��"9�D�2Je<}ux������@b�;"�)��|�Gs+·F[+p���Z���]��T����>3Ҵ\�.�.l��ly�J)��l��[��j
 ��@+�/�9��d���#	�0>��5g���^:Z��5o��o֠.�[�,��}#e��nZ���\L9�*���v�wHt���{m�r�ݪ�[��E��$�x٬�";�;9�\uw����,l�B�p/��ϫ��R�$	%H����X�@��Dǵ}�Y�?jL8<|��g�B���0qx.6;��,��ޱ,Ɇ?�)����C�g.�!���Z�Y#�F4i��%I�/]�垶_Q�,�Zd��6ٯځ7X�0ީ��63 =/�W��Į#j��jՠ� ]�
���Kpe�Y�t=J���1�q�Y�iM��8�Z��y���^�Zܬ	0���\N�֠���{���-�N��T�H�%m�'δt�f/&v��mNv�����ZU�wY{�E��,�bl����Ұ~��s5�zus'i�d��;�+c�4 %��P�\i�%p[,��+���޳\AE�	��EEِih�=�z�WmY#��r2�/{K(&?0�Zb��p�Z�� Y���nS[�]@X�jr��朚����W�9�f}���a>���%�8|��̚���o�B3E����h�B�F��������
����
��L&�}���	�%Jj�[h�f-�+_6O68ژ4`�aE�0�Z|Uʿ����<��6�� p7��z�>�R�4�)����������,_��>n����u�@�I���5�4�>!�z՘�~W�3�S}��4�0�+P��� ����#tZH�|=Y���+;_�	K]A�7���1r����x�Ӑ����2J�1;4�d�n��_��:C�弜�Z@:v�y0ZR��ݭ����8Ul�(�'o1 �&�gk����c�2�˰ޢ1_qi����`c��Ɍ��0�B|��=�'�m���.���bɚ�ؾ��P�à����>�<����+A<�*w���f�#lH�d]Q\U�<�����_����9�@4i��S���{���|�w�pb	��V.]�����6qu��
X�Gb�C�_����<�Һ*��\�+�^,����
�o�m|��5�y*vsV&	�?���	pc�'��Յ�֔MMGo-;��&��1yD�JE>Z��^A�B�O��c��i�EY�b.a����ǥ4�~�GHH*2����jf��%��u\��
o$��0:��Eu-ַ@؂�B!<-�Ĥ.Lz��w������w�n���!+�t�@�]������5O�=�n���2��;A,�~���ps8���v�j���c�J��J+�l�q�I�!Q��;�E������W�V��{�u�5�m��@�k�|>C����O���@:1+���s���>��!MMG� g��=>K_bci����Ў�w�&z*�)�T��r��+�ț�M�y�kO�D�ٗt��*���W~ӿ���qRD�$�)�a��[XX�ȭJ#�$9NN�i�wC����C�Z�j�!�j���`[�;̆��gu��NJԚ��^�ɧI��2 c�"�mT��A��������j-����wV��W0�7̫�u*>DeG����d�>��U���Z62�G����?\ԙ��j"��[}}�G3'���%BhI�%�_��M��k���[^K��B�¡2!W���bH]7�BǴK-��]P�ÅP>�B�#=��TRsM{D�m�$&A�f���p��Z���:�@��<b�/$�y�S�V�?Gl�����ji�E�`�\n�;�qj�
!W���@q⑿�@]�ٔ�9�;�3&+jy5]d����E��р
'g�CA���KQEg���㯶�Z�6CĨ�a����0r��2hg��Z\������+�rƗ!�ur���]5wob�_X� �@hM���:�>�L�V�q�Z�sue79��s��5���I]�FD��~o����`��ᾀ��D���+¢Sf~w;��7"�-�>�!�� �@��+����G��R���\& ��5��2!2Bf�Nb k0u��qkN�N�8J����F$�����]�|�@x�,{^<���1�¥��H���Z)S��>�W�Z���CU\��W}�����?G�8��ȼ���yưI g	�M��B�� ~w�,UkdO	��#'~�@��8/�f%��t��WwĆ&�W���$H���~x��ȈGx���nC^DpSC�8x��E�ٸ�¥�N��P������Q0%ߙ�|��BWW� 1�y,yA&���_�V6� ��\s�0x
��1�<l���s���$ ��Yl��+��������&��9�����>��v��I�$�
�����c���-���d��`�Y~h���+6�<I�9?��ޒ+�W<j}���3  	���s^�� a���SE��XM���E��f>qO	�
R�_� �MM�v9�^D�A}�	,w����C�n��+Z@5��o�TSy��x!<��'BU=��Q�Ro��SZ������4e	� ;k�ӼB[E.Հ�x�@�J�[��ؖ:�`���̮%�\g���*Q����F��E����![e���@���ơJ����Uܖ�br :Lt����ⱤB*�a��گ��%�Ѭ��L�Ա��Z&��2��9T0�f4�}�(��c�*2g�29�����>�v=f��%U��i�e�l�u%4��C�(�uXfN���}߫�">~�����ou=��+P��\]&G��G4��
.�tP
s�$�'�iv�حox���<C��M�x��1Q�<%�H�K���Ok����f�A�������ğ�;nY� �̔�Ԥ�g
����$�3]��S��?��\��[y���� {���L0mO�"Ҩ}!��8Ҩ�JH�+p�~����h&���[Ӟ�G~J㟣�#��uI/5%ػ��O�
��W�C���>��	�?�ṽSb$ږD��H��~םcV�:s��u�#�}��?�m5.�KÇm�C���sX������9n�~��q?��oV�U~o��{ؾ�b��A����_�]L��b�`�P�FFY� �m5�9��x�^�w�Bn�kt��Q�@�ʅדŎ6n��������jjI �f���SJ��l���m����!ڔ��'���:@��RO3�y?�!M}�?��}�)�� ���u?9� ����:cK���nN��7kP�:�ƔQ,k�.�<C9�_�ɉ����z���	��R�gbR�3Z��D�?�K���:#Z���"�� q�Cu��x�ܲFO�>�Uj��kO���m�Bi�����Dpa��O]̕_�ZV(�DϠqv�� c(���[Il���EC����F|S<��R6�)����9#��EQ�x�������w��f��P�p�}iS�ƅ������<�,WQ�DW�o�bB���'upyM�(��M�Eq�FGC�s� ��sG�n5s�9�k/n�؛C�#�Yc�Ӕ�G��
	� ���ۦ:�rU��X!��T��"�M3�!�<.L���՛|<��W���bs6EE.Yl_�����i�XJ*,�5��1*���K����f�	��9K��P"	M|��=�t���C$#	��0���K6��k��otD���N��(�Z=ƿ�|��ّ������5�G���+�����A2=��74�`�[&&��J��<����>�Wn��s.������^���VL�\0��q�S7%J�
�
�RR=�-�V1.F�c�{�pK4��/�'��n����u��dB���Jєh!E婟��7�'���F��(P���@龚<�$��EgͲ�n
c>��b�y��\=׉�[^����au�8F#>L�#}��Y����Z���Fc��S�,q��7ٿHJ��a?P���=�]�Z
o?+�l��%g|��F����
�#x]�'�����Ol�t��WG �#_�?��)Ձw��RM��?dIs9|[-��'צX�8<�dl����Q|�xC�X���t��V��j��0e�4ObE��+��j ��}�)w�j_�0`)4AcV{�p+���㣹��.%:��R��¤J��Hz��U��b���_R�c:�(p�pW�1e
	̀��0p�M,F�0�)5=JFpw�d
��sGI}gͭ���tw|�y�$Y�T��Z�i�xĀn����ȗ]��L��K���O�Za��� )�����:��SF�������U1�����Qݿ�eF��[�10gj� =��Y���)�B�QƜ���sش�����Uf`je{O��L�|�Yܟ�n���U$D�N�>E\�7Q�]�6z��F�3b	�3�\��Y*Ub,C��!n��1xo�Ͻ~�N�%����h�<(H�+�U��vB�� fi��&�FA+�V��
�kU�Ň��e��s:�,��Ւ�+�~\���r�����j_�a K��Y��g5�`%N?YZ�gn�3�Hʑa��_Ց���:��}k�!<*�f���넌�.��~�}��J�jfgB1O��aeq���r���<�^���$�"�U�?�� g�l���@=E~�ņ��y��%��V{��h��7����r �bL�I ���pSDD^�����`v~�ْ�JG� �m������SĔ�����v�`�ʇ���1�z�C�|)�B�Y���j���t䶓�s;l�&��w��>[k{�6*C}lF�#ؼ7CTy\��[n��l.�!e|m�[[��v�r"�o�M{y[���K�� XU���?�sR�����$⯘Һ����uP�/�W91�(k�F���J�W�hR�-��ռ��G��G���3��(��P~alR�d�2!T��_���\�ϩ���z��!BaZ`��5�e���K��$5�|���k�{����=���x���rB�;'߉M�e�W6�f��%n}�YF�pab^�'���sIL�|�.7�x��Jpb*:.�/���|F>Oĩ�����>�IƲ�T��'���~ǻ�}��K%�	����F����)!m�vo����K�B8,Qv^��8ns�_����	7�wl���6���������ڱ"��$�oh��xJ�ꛜE�S���p�.�(����kl�4�I�D�A%-'A,�����rHNW�l��3�@�y�#���0��)��[�2Ⓥ�HŤ���r���OIe���]���^�'�r�ދ��u��]�D�����~�	Ie	�;����g]0u��"ʦ��UsI,Ϩ,�MtC�So�S8W����*p�ơk����p�|B���@ ��FSaП�"!���b��Q���D<��`=�s�����"*i`Tːg4�9�Ɓ���R�3��`0	�s$n��b37/DyV#(2~"Z�������^���O� ���䇭A��X �U�T&Ĭ�����NϨ�Q�r|��S�Ȩf�c��M��հ��XU����h�c�ڊR�B��s�p�uC�����~������ǔ�K�����f��g���]d�*?����X��fYa����j�L�\&����R��ߡ-[`z� ͉���n���-�K��QP��!0��Ͼ(�'�&�v{�~1w.v{�G��%�Xs�w=��q��+�7.�8vɫv�8PF�Pk�=�Gr[�J~ZÎ�V�Mv����>
� ��O��.w��	����O�<ڧ�u�������q`_�o�v�C��'�(G����f��C�5���;�W�)���4�><�K�b�"�םFi�LOd�� w����Ņ�`|o�5���q�i�N˾Ĵ�:fp�s��-o��fV�{ܥ9?ԓ�o�l��3���⳷;�VZj���D�5�D�u3��.�O�@E�Z������k-'����2d�&���Aʮ�e�Z@Ÿu�V� ߕ!��0�WS9<(�y��~\�1Y,V��b8�ic�v_I9��o�NAQA�$��pC�5*%/%o�t(�9�,�u4��b�s��f��7|���5`'9�������x��;c�S+ �R��091*?�����I�����!� � Z7E�h���HEE�ң���uX�S�R�w4N�n�S��ui� >�%qq{�Cֲ�F�t�����xr޴vi��mꇪ�= ��?�ͻ�%�F�HQ�;�Y����sz� {=�'`+P�_�a�|MiG�Í�,�!�V�����H"ܠ�~�<F�4�}�HSG-�!�U���Zu��ŖbV�y��qv�v�y��9�u����@��s��|[�e��=��/i� ���k���x�c�2����Է�g��m-qWݳ��k�e��@�d(}S=$��M^r�=��J)�]j'3���S�z�U���
�>/�NmaI�8��W�e�`��f��?��|�^�'�Dj���iϏC����Em'h@ױu�r,qq�����\�%;��̒�{�GU�X`e�׾�7G�@W{g-�S��E�r�ڃ3�u�(j��%��+&�1�E n��+��z 5h�t��΀�{�jOMM�����a �����{�0�YC�U���) ,&���8�SW�¸�\����*��N4��Gi���=�n�����`�?ҡ�
����?v�e��-Ŀ�1���[�y�PZ-�F��O
p�? 6�Id�����euz� w�����U�9����L1������Hh�LNb0�b��)nؼ��|�Z����v�����2+U)�q�n#5<g�郕���栃�1B�[�,3G�tb���z��d���+��W��>�f�U����`�p]J�EmK+��I���G�L���A�w_���P@��}D\���j�3��_�h�9c�
ه`R[|N�x�Y�a��ϫ�;)�SV?�SZG����D�")^��3�2�����Y\V�I����*��b�ρ ����5���
�2,�i��ۖ��lgs���z�;�?N�Ћvf�W`#�*&�#o�1 =ҳ��)@�3gN��� EZRk�Tǡg2ȶ,	8��Qϴ����'|	�O���1�q0�/��}!d���˫�`d�n*��$`p�ܰ��<�y�3,uX\���~4�.����Od��Z?�:���Z�c^s�q�mR#1�k��P��-����1���t��r�wy;����e�c�W���)i�:�F<�������Lk,EU���%'���0��Y_���8XJ8�؏vI���"Ɇ�T*��G[�	A���t���"m��EH�|T*���n�'/�$�@7(8�U��������Fu�5�46%��s��Z�t]��O��cR�J��� �k�M���W����^�+8>ԫs���ϸ$}��>�H��c�s��ݧ���?��Z�o�q�K��q	����jÍ��"24�� ������W�P+����衸�­c�O�k�w��˺�'���pb�f�����������@�~���:��Ojt|����F�����~ ie�\Ժ+C��}��P�����5�	i����0��Vx��KqS�8�H̗�)��PGlLtz����b4u�|c_���t�L�&��p�A2��D)@��d��8��`Ō�:s-A�!���o�
����*r�{r��~��X�}��d���<�����R��Z�(vS�q8̯IO� 7 ��Kj&⎔����%8=�����k�G��\/�L�Wkj}�.1�	6�U�Q��]��ot���	����	��c�|��E��w��T#�����$��������NX@��Ӿ(t���9����6�<��2P&JӠ�����۰MR�M��fy�pʽً��i��w#">�.CVܔ�'���g'����Zi�AXfZ9���E�[ �*	�+Ia'�侷%��~��eB��~����CC��<	U]��0�/�xa�u�r.I��d���W6#�����]b���*3�t${��/��"�қ4E̰�
;u�.Q�#L�$����ѻ��>���ָ���:�!�$�5�Ͻ��C81�J._���0@���YK��*�k��I��+���n<_�z�j�x���L����7lN�}y�:��Ś|��������F�b�L:v��^���@į�g�I@�s"p�6u�c���j\|sC��Ќ5n���3VT��#c�����+`��:��:���R͞�t�+Q�-������!���y��{j3J+sB�k)~�_hz��V��\j�T_�П�4)����Q,ba��8�s��1o�-躆��\����,C���߂F�2WT��N:�-e��ib�;�8��lE/rm�;?`�z��]����/=��s�ϖy����RE�x��)�,��Sn�{����Ԑ?1����Lp"+�-��g��{���JÅ���|�{��T��4YT{t}���Ӳ����g�Z���G_M��L�Vv�k,���c���k.�� �-���$ro�=�~O�h�`v�G�y�D�X~��9�,����_i���gq�� ��Ӑ��3�z|�X�ȅ�D���pY˖�����ɦw6Ѣ�q�o�爼@נZ!χh�w�3c���f֠X4j��&w[�Mk��B,4�K$����KBn�8�P����!��J��]ɫ��8s=V�3y�X�œ(�}�����S2欶��Z�)4��!����˴ƾ��Kg;Ɩ�"d�	���D@C\�@aX.I�Gi�f%����u=�7*�'{ʚ�>�0g���	�뼾Y+��r���rH�9�Q!:�M���ݱ�t=^�G�V��
��óo�;���z����������uWId`n(����z�p\��Mj%��P���'f�X��ƑX��V�G�X��f�9dг[UO-w��~������z

��-(͞��8c���Z%���.�e7/X�4F��ԉ�8�B�����UR �y1���v,�
��i�j��4���Ki0�����ڴu��q�� ���}�S�g|텔�#U�7?o��.�~��CA(+�G�4�M�}m/������쌩�I��dgوcz`�W�J�Gms���������M'��"�4/�S�]���Q.Y�M'���&w��������.��� ���txxa
tg2��sV��Si���-��؈��G	 ���]O�����;�{.b��)��-�ƾ����n�\Ԭ:���B��2���yNZ�	���PC؆U_5�cg˅��2���wOc�����pí[Dv,�[G/ބ�Ā4M�!������_�R�k�ߟ�p��r?6Z���cj���'��R���Ie|
yD���l���f3�-]���-:�q�'s:c�?vX���7Q'y:�;&�n���9��r]֋��q�u�W���u�<���Iz)�Gp��<�E
c����S���Mg���fG��t���/�O��/��b����8�tA�X>͒�?Ɇ|���FJ����B�	���s�O�?�v�.QTK��RS��z��~�5��8ʝ�� 8�vi�4��3��G@#��D8Ѱ��W�$m�"\��{�r��1>j���I�C���N�9W��I�s��#����"��u���	F�s����_�2��A~�-�3�ǘͥ���_�>�5M�D˩���`ŋ����ȶHa;D�^o���e#./X�F-�����O��K �_HR��tx�[A���Ea�|8��]K����"N��m���oJݦv>{.f�42�Hk+����Wu�ܗV��pr>>Ut�!��s�>�F����i,���P��5�����8��l[��%���t ��1����ց�͔HX�Q�h+��=.��i�>�M��mg J�< �%�bi��O��S�0��k��u��SQi�D�&�}�G��WNN�S�
�>7;AYݎ��:�gW]	�)z��h�b��f%�FZ^�ꐙ����v4;J�4�e�Y|a��st�o��<���⠶˨A'���s2I`{�T"��D\�p�`|!�Fa�!gf�7�=d��ʗI��t�q�������b�'����U�\��7�\N��$�v����f����-�:?�[�ە���p&܏"���!�f�$u�^2�DyAz�-�ߚ�t���?v�Vk��z1�/�Uva�(b�3%���8 -3+�+��9�<T�Q\<	��8j�����R'��� �����X`Q�x�v�T�s��WK��k����F0���Q��$�lD����^Yϸ�L	2�=e�|��4BZ���e����J#��ӹ����輻IV{O�Az�c�xΒ�9Qd
4F�����:;�����7�}�� �U�zz,f�iM��\���Y������fr��[����%ԉ��F��嫥d�����1+3�igY�?��.y�i�!y��,ڈD0j�'=� ��#<��àQK�҆Ꮻ:F���FM�2�l:��#�DK�K5�z&�3g;Nr����3�h仁�����ա}�On\�qn2%K9-��r\���`�I:���A�Ђvoy��p�*��� 5��JI�<r\����.읱�
k8����5�w�c<<K&��]���n4�`9b_ ^9Ox��2)�n�Rx�|<Mo�����N-�]�L?2k�G.,�y+��]�J{��Z��զ-F톈���Ux���HJ�F����wɅ����\��&b���^ؘ��䯱��!� k�	��U����9�N�B����d��A�'�0	��ާ+���3���up=������;���N�"��X%*皶s�f��:�(3Uz�,�U�+�9׏��M໓+��R��^�]���lƳ�qc6��i����o��B�8����.��2l*M�MGg[���3F�t���[�ߝ�fKks�u\��;�A�Xj�2^�>k�u��% M��T�arEb��������*0�ݘ�oR�\M������צf�m��B�u�n��A�3=E�|,��(x�@�Z/�7���5T��-~�t>\+�0ڋ��+'غ6)���ե"��$�Xx-a�g���ݏWj
(��{8�&�r��(����7V���S����:�Tء<,��A<wf�{7Ӄ�l��A'�ˁ�Zm�z#�uD�;}�ut���Ҩ+lmi�lѸ 8�$�&��$0y�c%b#���'�J�a]@x7� Y�%��Ĕ�e�Ou@ͅm
(+���V:���w�
�_����I���<�:��FV y��ڻ������B�=���s������?/�8�
��^��þ�G�����~s�іVq�;��ϩ��p
g(�x��}�~��%w�. ċ�ؽGC*Z��8�%��Y����a�E���گ�����ί�oI}��Pk�,�\a,=O�޼���f���c��ظڟO<Z�9��헙-a
�Ur��W?��p��sJ�[E]�Z�����1\1SqZ�	wM��Ӕ��-�!$�0�F�F=�)�Я�ەD^�R�>J�:z.o��hC�.}����Z5Ȩ��)o�Q���+0.�4�>�� �%TFge�W�꾙��BC�*��ۭ�)\�|�!5�)�q��`�,ˑ�K,�������.��}�x� ��:Q�dh�vV�ưY�[�W��Wt�V�+7���������D&�jyE��-ԂF�SAK	qO�|}Tz��oe��$4�<�7(f"?d$+���yU;��i8c�决�ʦu��N�ƎKp��sJ~Qo�k��H�;��T�k���?��]|��=�~yL�-؈��(�rTb�:�I &\-H��?��d�������<���������鳵��{��
Zq4�� �s�%N�D#>�Z�@S�+l�t��^��ޗT�Gت���`mWg�7�)�#�p1����-u$���"�1@.�5���W�M�c!\/h*�����H�����;HM��)y�(&/�������Bb��ö߅��E%�N��~��2���#�* ��!��3K#O��T�� ���9�n��l��������<�K� R����w�/�W�jow�y�E*e	�����HF�3H�A\H<�RDg�"������D���c�8`z&ة���/�����o�����I\�$^�)7�e^�~��Nt��w)V�|��֬�x���L�ڂ�]���i>r _��
�T>�?�R��%F�>�k9c@��m�q��x)[��ʑH�̼QD��zzj{�|�u�Cc1k��vjF��A`��t#��E�<&n9%U�CYG3<͎�}���-)�j3���<�Q%S���We��S���Jʎa�[��ME�N�p�t	�{�+v6L	�o{K1�_�����,� C�/��|�>M�4�3����z�\��Y>�g�����5�}�rDЕ�KA�P�����2`�pc#�zB�C��R�
E.���F�J�����޼�h�N�9�q����K��$)���=V����Rjs����I��-��7�n��{���;�9�z��H��pc���$�!7f�$z1���<h�)BVTZ����'!M;v3�>�]	���c�^U�*l扫{�!��/G����z0L��*��Ȳ��	0�YXc���S��|��~�M��d%����%9U�k��ƉT�J!/xnt�+�v�Q2��	�ӹ�V��mt<XEH�$(�Y�"7���6�n�u�;-ő�1.83�K�(���߱�i�>��$@c�_St����I�Z��j�	��զ��q��kW��ǡ5t�;�7�� '����Q��z���C�������/��Z��F�
�J�&/���Ͷ��O�}���B���3�:�'+�� �O���E!!F^f�5�7���b|��-C,Gw��sW��m��T�ծ�X�A�TT�9������?0��%�3IV~�W�l_�i�����a��1�`7�\�M��*~�C�B�n��k�m#�+����g&�T�V,��+U-`�anLm3��f$���@{�����Z�9X��1���k[M�b�x���_�E�%3?>klS�����~�:t�x*}�,�c����*8tI��>Ne3=�	�s�uxdACwF�+N6Bfr��G� 5Ep�^W��,��vN��.�ڬ��(�Ů�tT���Y��z醛N�P�݌8%`pz97�/B�V�p�c�c����%�b�	�"�Ǥ�����%>_<�����{j���¾̒��(2�q�|=��B��P��o)}�	N�o����2���_�Ѻ�L,��B����x��ٰՖ\1c��!�p����S^[�XJ�N���t�M��� �1��M��(�A*F��]f�Ĥm��Z��%$�r􅢭�Y�Prm����Tf���8���gX�WZ���xgD{�TY���Q|�=�=r�}�\�v�1�/7�x?.�������;@-چf�ݦ���X�q3R��Mp���2,Rls�����4�]L�-��̐�`:����i�L��f0K���3���%�D	��2� � \ѨŤ���t����(����p�F~��V�W�+p��X)�����*r��ʉ8T<Jlb�R�P�JjA�y߫dۇ9�R_[B�� j��4��3M<�Xu�%E� �)�j�~d���M��ω������1I�<���1�»&:���!6 XtZ�=Gʋ��z`������V"��k6 (�7T��
��g[k�j8��M{�%�:U��i�������-x�\ �y�c���*8�,��É=�5R�Z�c$��Gqla�GD?��P�n6ލ� ���KP�\A%�
�M��<����\�)�.]�6S&� �'�]�咇8r9��ɐ�D�X������y�ɱ�Ug�~|5f�nQ�[�g�U�y	��?� AHEs_c��zy���9���9O��J�kR���D�E#Z�Ho�p.�AJ��HH�?4\����^~�Qą9@��S�Ϗ�^��2�_�!�Q\��F��<2��-Ņ/�wj`��7����4|�ȼ
���r�6�H'���	Q�(h�rV�@�P4J�r��<�
��$��j�1���Ԩ���x����<D/��Evв���Cpi�����8G�>�jOX�����-u��"uwo��i�M�����w��g�U��]b���Lty^E�F���W���l�V2̭�Ҟ����ҧ�څc}�1��/<S���?� �Ѱ���.�+<���5�'W}�~�RA�Q��in9!��P9B�n	�l����l �z�/2(VI����Ŧ�t[��z�� Շ3o�ig��bͲ�Yc����wcφDo-���D�ސ%(�+�F\�
Y)�l�!�]� ��k�(�Q��!�ZC*>�8��்�=$�rͼ�~M
����׉x�}r�#�!I�JV����D��5x�DE��>��� �wؾM�'��Ȩ�=���k_�����V]��A���&#�!X�G{�+��*������(�D�Vq�F�����a�zBNzE��xZ���1�6�荚mpS:�~��:��ȕLJ4�;�����'l4H�gַ����ȫx����-E;��OK��E%�z��Ȉ���]�n��M|���W�uM"0bD[�H�����v��֎��[�]h�,��5�&����%rݒ<���O9d��l|ڴb���f.��yK�	��ڠ��=x:?(�r�Ks�<�}�T���~�-ƕ�䅵h�{h��:u�����鷻=�����+����������v��P7[p�R}8����C[i�}�I^`sߊ�!��&��`[ ��4N@+ʂ����Ej!�y�Jf����/vtQe$�m�M�3Ϙ�b�mGϦ>��4rM�ߝn�!izޑ�ź��b?w�A�߀�Cx.�@�OE���e�Vz
b|8G@�%����kF@I|�X�T�Tp=�C��B����B+_,��#�|*�;�C��@�Vyt;v�q_�����Dg�q�U�,4�2:׿���~��`TF�8[F1ُ7���[����3�Ś�Y�4���j�{��ra�"]ô☷��o��|��.�mGG�{����u8��G�`^<_�+�\��
ޜ�����(�8�\��Ы�\��<���{��Q����_3*�%��s����}��B��"8�ݴ3�dtqX����I8ķ��i������ !b�L�b-=%��D��mV�w4u��6���{����a:�!� �Sˤ0�]�����f �L�mH�Гk}�7Bj��~&��D�&>�@�d����-7(�rՕT"�,"]r|��f4�F��Ft�_��lAP�4�V���x�Y���ۘG�[|�m�	���e+���2��G�J6}J�^j�g���|�" b�Y��u�Gfx`��{�[3߇��LU�����Ⱥ>�<�7.�s�桅��C��v1�0�\��9���U�2��A�*3�|�ܷ�%W֡=�%�����M�ر�Ź��Va�-@ǔ�b����S%�6��obU�n��{&�T��CJ���v��np�Q����9IN(�+���U?e�^����2l{�
��Y�1�k��D����� ��b?���~�.��pÃ�����̡5b�e�Q�`H�n#5^�?{!�YrVs+:C��!lFȊ��\�,,�V����֢�6#}�i�ne̿�S�)��n��ۇ|0z��z�x3�
,V�-dwf��2+=߈B;��ۉ�'��IK*	��̗3�DmK��V4w����iˍ��V�@S�L��ƒa�]{'	?��s<��Xd�R����WqB�2�Eʈ���.8a��c'��-�jo�-Si��M3��ʕ8[@�7�ڹ�V1��.u6e@�?,\M�m��9��ZW筢q�ʾk:��I6��m�.���e ,L'�&��ė��j.�H�;��|��:�`kv��tܮ9���5SK���nr&���� ($X몹�	�3s�	�L�&�zF*m~^�c۷�@xzS$��t��d�h����,��_4x�a\%���ot��AȎ��� ��Εg��$/_}���g���s-�vc*S�s��o�Y-mb���&v����i�S�QX�N�ߝ�KNO�E�
9���%�� ��٧���lkIa�l&��rS�4G����W��("��uaA�d��$c+�c����[�BhT�a[����G.$���:y��l��k��?+�\���9=��Wѥ?�P��rMCh���^���$m�p:N�������iY���s�#����s����׃#��N�q��~ƞ�14/��I�*2��r�{z]�v�B��۵ts�r>�S�v�_�����Y�Te�V�Dn8�h�>V⽒K��G?�|Q���h�9�]�v��F�3�F�:.��ݪ����+X����ݹ1��?^񉒄�A&;�۹�8z�p05!]���ϓ�/P:s.�Z�n��ϖ��w�C�n^2���"z�����������#MG�_@�i�e�Т�HMQ"v�.���I���~b}_qW�rs���Zo���v���ݬ
��Cd{ܓ= �3ؗ0@͸��EN`7}����2!Dg�-��:�����6y�yG���IUx��F�ȑ�Aխ��"�Y�	�L�o�D�F�>azTo�G�����_m�^<Ŷ|7��I�z�H��NƊU�S�ID��g�pcM��<ls(u��\�	Ui7�2����A��p�3&�ъ���Z�Y�F�2�P��vA0�)�?�q���� b����lI(�K��Zjg��uߨ�|{=�"zz�GOȭ/6ӳ:�s���D&��G5u�E�9�=7̷�B��>�e"�TJ�O={R����Y��}\p� Ғ�3Z-=v�L�%��Ko����/P�l�QQ4�TJ�ޤ���t͝mHY�ˠ�B;F:�}H�~qizi�%�B�S:,�O{.+���]�ě�������Uש��������y�@`�v��շ���&
MT�ڕb����2�S#��B@E�%�4ei��D�s��K���Ɣ�0�ңq�u���Ny��Bx$X�$M{�ފ�e���v6M�i����>�г@�a�am�4��62A;$��u���{+��T�v���HD�y�Q�0� H��vs��[~�H1�zK&�4{v4mRt�=N��!+Y�c�l��}ɏ��ŪH��s������б�^غ�2t�QY���H%��?D�p���
4����J՘�Dt� �r�,�y��s��ɖ��
�c`�4��=r]P�7/0��ld�$��Q4ŚÚKq���-o�Xm�Խ�z!����S�������Z��7+�Ԏ�g�+tM8n�T�	�$�sa�j0�v��T�!v� S����=�Ѹ��tG%�o����Of� �W���>��)פ�9au��tK�o{S�Y�C�GH�{EQ�G����`�J-���f���I��"%��3�a�z�G���,2cb�M��|}M�B3<��#j��\p�{"T9��_t?k���D���w��W? �Ԉg'RJ�f(�E�$x������!��;��o�6��¼|�m��
Y
�q�3�*͂sso�ud@��k�n<�����u*?8�nXϳj�)g3Ȭ8�򬞲���b�O�B��b�8&%������Ċ�7���0��4VZW��0FI.`ţ���:�PA�@�b�����/�r�-��w� ��i�<���3��I��+�ly����T�A�4�XCSl@�Y��8_{`�pu�c$!oԵ�՟�-]��t�Nh�MKE�c���6k�q��K��ĭC��'�l`�����i%Kk��׭���c�������"�`�c
�-@/�%gLP��a>��oTB��lK�4��9�i��<w1f3��w����zX��3 .�*�$�z�!>�ߟ�e�qu�&�� 4rE�U���>������_?�RY<<!�X't��v�i��Q��t;/0���f{8q(2/�Ќ~�b���"l+�QdY:�"/�<�̇�`������F�e�"�L��P���5�P��5�{�� �c=����G�`�n��d��ߊr�O֗�\�r�"a�]�W��3��s\��[kÀz���"�צ���=��it266�3�$���*a�+�'+/jG�5K#������
#@�H��汃
f�j0�У�@e"�P�%5Z�F/�F������@�����	�M̔�IG1c���e��"1�DY��coSEC|���ө��2S'+!tU�',�n;��ZVvW����<���0�#����;PNb8��2��faM>�Ṕ:��"�`��q�߆�qV|�G���
�,����r2��;~U�}+'�� ��\EC�,� À�*��%�縖�d����<O9�"�A��u�sx7��9��7C��7�p�j"�KbQ=OY�d���.�	밎�߄!I�q���A�c}��+�A�l���P�%g5c�/N{�u4��}g!��#Z~�W���U Z�ٸ����E>�,Q\����t$�tя�u`�.g����qN����bվ��z'/�M�c��d��3*^ޒ������r�!wk;�64ck΅-�/2B�Q?��)�/ܹgL�p�0O�Ɨ|g��#�Oj�̐�,֎{�ϗ�yzmj�c/gW���	��eh΋yΟ�6lS�ǢGYWr3�y+���
��Λ3�M�7���;h�d݀~ VJ��>���AB;���h]�P�m`7�v���d�c;����Y���hǹN�e��o۔D�:�A����SoBǵ#f-��8F6�G��r�	�5o�딁:#
~- ��Jͣ�6��m8�s���N9r�B=��$�C��H��u��0�
��K��K�7�`
ɮ�:Q������&~Y!��J.�&D743\��vm�QB��8��*f/_��Eۄj��L3���ۈ�ŴE�'v�|5�������e�ys)ͭx�;������W��� zo�t�~#X�L�jy�~�׈��`v̕c��p�lS�a�G�Y��v��s�����z�mC-"Qε�p��G�I�1��Y%��P��.��Uh�	@��
�XZ,h��B+�z�yA�#AUH������4�*�X΍~�K�ў4x�'Z����5[��!M��g0�B���+T����6�	2&'r("�(�y�Qj��<T��7�>`��u��IA-���ƽ�{HcNt0�H=qn �N=b�'B�-v>.�đ˚�F���������>X��
�vK���s��l���-���g��t���b'V�2�̖߳�e����s]����uQ�	�E8Ԙ�	��[�=P��X��xW�u��ȳ�R�7��k��߽T���\n6�[�� 㻵yD�</�cy�'w�;v ���&8�Qg��e��2-�"E6�QbM���6��V,+�6F���9!K�[���UoH�FF�@/w�;E��^��<B�.=�b�g���{��x�~("��w�ܩ^�	�w��	��,��Pʱ�	�ub"Tq��j�Ҩ"ف�5D�p�H��	!i����X�eݼ�O�A�j�=2�+�U��&��r��z��]Ж�C�"!�g��6 /��z��P���9�H����?��/�2�f���@�
s�OC�c�\}�brFY�E��(&���U����=c߲<�%�M��lJ
�륪�5G�
U-�TPoq��P4Mw��g��B��x�$?��}�$ʉ�|D�l���S�����f�ac;�9k\M/����w;?Lz��u��vm���!Q���]�˧�+*����U�D�P�ci�(4�߾c�Q��(�|�Sȡ��>z�Zc̮2<�]�+K:b-�_|�>�̎d>G�re�"�:G��}��b�K��Cz�b����r��O�Q���oE��h���Oa�S�u5K+!d�z�{}	�'�BNi��`$�ܽ�ߊ����F�s�_TPȀ�$�ƻ4iσ�ť���h��S�5nC�}�o�-ɧ��*���w�0hVw�D%`��C �w����e���u�!��:�4[\7��p�3���KF�=�Pt��9�W�WO-�E�E[���h@��QǤ�?���3<�v̛U+��Y�!вh�x���F� Q��d�"�٢�\*����ܦ~E�2����s�Q�����p�Ũ�0c,/Ւ�k���w����N+t��NQ��A�
��d���������:~q�x&K�����ֽc#�`��1���+�����_�kA|�5��3�uIs��z=�� p!w���fը����d���=s�H�ݸ�v�ۑ�yk��z� �l�x	��{r��cz�13gZ5a!�>DЯ���FHPG�²�sr��}}]�^Ծ$X��@�Ah:"�Ġj��{�ڑ�k`��9��P�yq��E���npR��%"IG+S�˄�N�M}�O�0��aBPr^�p�V@���( !��Uh�s�F���!����N��r[�,�r��X��V�<r�(�9���2+����-G��B]�ӛ�|���� Fm�k��[�/jIֺ�S9�����U�Mj
>B���рBX5�XL�(ƞ����Go>6�w0%.�b���aE[FQ������瑀
�q��+�	f`�8v��� I���dq�O[��*�L�U��o+�:�T,��{����e�1,�Ҵ�$"a�n_3�[\VȪ�Z�&2d�.j��Qv]E��n�F@,���|,E�!��Gw� �����D�A�d6n\���A�P/Qby�Ғ���e9<PSK�پ�
���<�`�z��<Ү���w߯���l�|%V��8O�.��Hv�k2�[Y9B��:m��V�������������ظ����!�b�a�ۆd��Y��oXK��x�����l��mA�%,�#�k�Hec��垅>�k��ނc���v$V�od}��i��M�G�O�d�7+Jk�/>��{À���������:]�9o�u�j����ɹ�N~R�2E��3���)�h�+�¾_1�W/ XZT�K�hCb�3.o����c�#�j(��3���9<R��e�e)}}e�Rcl� ��0���a�j�C}�9btM��C+r��jwį��]r�Yր �� �����	�:8�yup�v�~�vg�5=�v`�����}g�Uj�����/�S 9B����0�+ 9_2�����m-4�+%�I�0�g,F�єr��\R�sb�Y��ɨ���{��=��8ak9��j�޵�T-���Rrm��u;DR��逽�h���}�\�}��:��ĄvV?��D1�=����r��:�2�D!f��?�sK<!���1�����?���s|\3�i��?��phB����2Q�0�m��C�
�)e�T�J;ez�i��N�w��\"�zS�,��̧���Ʈ�6�p����pK�V]���s M������h�q���0��pķ�,c�#�jM�w-S� ������GYh���Aۛ��1�������gN���EV�_�Ά���R�<��ݳihgd��9�y��1Q+̀췉�A �ck�WN�.��2{J��28�Xwr����$z��<�)�G������k�	2����Ev�8�rn�ݵ�~3�I��I���r&��P~�_�'�>�ɠ���<�X���z��`���}ABr�=sɺ�5��`�������.3�jǔ�(�`\�Q��G@ ��{�'n�\B��ʓ"�rh`��l�{����"�%�U!θ�f-K�jq�v���'I��������M�ELf7��׵�P�ݠ�c�l�����[�k��W�T0���eiù.W0i��K,ٌ���%��Zz�<�2��hC��J�#)�o怒�ת�H	&r��#-�ߋ"���4n�5��#�ܵ�9��za��iloS7���fr��.�V<���0~E��p��j?�������>)�[�e����Z�ڃfzG,�K�>1wˀ�P#y^�͒��+[\�VE"p����}�VWX`����0�P�ْ��4B�o'�°����p� =u���낆&�u�h�z�/���\'�r[���H�B_��s�7��@�_M�E�{=�s�X���M���i��Y��D�'���5�GT- V�ogH�f�a��cR�PLr�m1�n��#G�?�T�u�=�gv�O��B��}�ұUs+Pfu�dUw7~}��(�a��z�ifg�&���+0��Y�ϵ���	�Қ���sR�B��"���s	��4�IM���󈓾|؍�����E�	&{D�-g��~���7���v��� ��|b��l��U��k��)+��'�Y����>�ͯ���h�5�
C ��%�R�U��|��2�#\n1�`�"G4�S~�D��� ݚax�L�^�Ώ�9#���|z�Y1[�L�s]`���{BIC���9B��5���HDۼ�&���YE����>�D#���L0�"������ݚ���qK`�RF�)�6��ތ�5��� �;s�Wr��#Ϥ\�[u�q�V��M�y�@�%kΟ��
ћ�8�� ,w�|���I�	����z��_��ƒ�0�dZ��]���5r%]����l�@��h�t��W�*�\�Tc�tNH�G�����J��q�J<���-�E��,Tp?aÿ�q���lQ���m��b���4�����#�+�%^��L�Ȉ=��}T	��o���Rl���Tʙ=�l�]�D�'$#�٬|N�9|�Ҳ��K��$y�U�/A �35�&�6?��@�-BP�$=��8�DVH�eٴ���`LW��:wX�h�W�[YO<�R���<[";��|XՌ֚�y�`��o~�,zc��=�ߞ(�����!hm#��w��"���q>"3b�D9�9C8I�p��O�]�o_�+KLU<<׾�c�Wxb��,������6�^��QPH��ɧ�������B���`�j5�i[Ln��R�ڹR!~Y�Az���vxa)&|8n���[M;>���W��Y�X��+�YE��$s0m1�~f"L<�	ؐ9?"��p{���پ��0��BJ2��N �)nvu����G�0�0:�)E�¨�0p�ԋ�o�Y�ڭ�x��+7ɯ�2uDA�ˠZ8,SV��u���خ�L.6�Y����8~�0�X�=�M��e��(zx۱L��������?]�n�Z��傤�;�U��ǩ�2�_7Շ���f�� �  l/�F���d�mY�y�v��=���/��f���s�5~g��������i_�A��1h���$Nu�h<�[�|tzd.���_�aʔ&�O�@_���rh�����)(�m�� Euy�I��Y�J���h��"bB���;Gq�L� ��elٯ��+:e���$:P�L[��u���_�R� �����Os���f=���L+��Qu�h�Y���[��t%���|�����_=�����tQ)�^<�I���=);Ă7z�Ft+caأG�C��33��,iN�rKˁ< s mș�
�W!6�۸A�?y^z�I�5�'4�A�G�4{u͝���1����
�t�m��pK�  �	��.wI)M��Zmز��X�+��˔���׀u���v�!t"�n���A��XF��z3�د����ԓ�d�\�Ir.��;3�2j��qbŸ���J�J>�:Õ����8���ޑc��^GAZe�1��1GXcY��u"bI	C
旮�B�]6�D�W�nN���g�_u�	�u��R���,l�Ppp��F
t�Ƴ�7l���C�`/�GI���58�<�f���K�)-��L��ɟ�V2�h�R���6Se0�)���DS����o��{J��+j� �oȞ�y������2�3�=�N�'������~�L�B�%���=�B�X�ޯ<�o̺�"��<�Yr�fwyᇎ�5��_iCx��bS��X����M�̍\^��yXV�@�m�u����T��% Lb�ʱ)jؑ�h$17�r�=���j���O&�WNu��'ĺ�8�	(�a�o�%����2�%r�!Q2`��]/U*l�V���?.R��]�3l_��x������TR҇��""��73̞/,+LHh����#vj	�orh�9�.���4OT0���g��!��Kɇ�c#�ĺ���3�tR��^D"?�T��_�=�s(�p�P��2�K���ѓ�\,�03�E��g�0�LN��`�5<L0kq���|� ���\�LR�	d�~�2��g��Otq��CU��X�u���K�;=h,aCc�$�������O3�ߣr�IQDyf�,����2�vG�ڏIk�i<��,($I���OD�7ݾ��QK.�k|xn��O��ո�� ��z5��~z�Gq�Z�5>�0�Z���G�xdcW�}�/�\o\��m�^����.��0v�秤�	��r��B9f��!��'.E�־,p4�U���U6*�ծ%aX�n]����횤��.:ٯ��A�{M������w��(v��d��+x������ e+�}��YS[�D�K-ΞL�B�VL��x/?Q���xw)�ܾ����������ٞHgs�>{Ք�����c .rMvd&�p���:5�(_���V}�w�Ip��j������@j-�
�ͫu����D| �)_�{:0�M�%k��ɐ�������I/�q�`�Uf��=2z$>�u*R�eF�o5��� �!4�BC�� {��Ѕ�p�v�n���j�s),//��xu�#��iTkG
z����H[n3�Yt�T��@QSV��r�~Q��PK�/�&�V �(��Z��q��wk��[N�}�z����%=�e~C#�n*��N�E�N��d+�MB19+��Y`����!R���ѥT�TJ���r�F��:ߠ��۔�A������� �N$�*C�����H
&�poa��g����X�ި��d_-�Ԙ�u����1�z>6�yM����F��9_/v7/IcC{D�|�繼v�?ab����D6��&�e�3�q�~�=����|��h�C�Ԛ	^�!ճ��N��0$.�Ɣ}`�}��Er�D���8���X�~�c��W��#�x{k}ι�k��ew�-[6H��<�$o&���ٻ��;����V$v���Z�ݸP�0}z*D����?1#��]K���w���4Ў%Od�e�Ӄ~h� x�^�����wu\/�~	��!E֢b��6���X��I����8H��OA�Ϙ�_�a�F��H�����U�i�3���T�EB�uO���:T08@y����8���Uz�i�\��?6;������,|�K�z�R;m�{�M3��1�R�vE�-�Ɓ�r�Y�&f��S��w�^�ik�����'3?��Gr�nI�'�9����Զ���� *��d� G��{���২�J�&��ob� ���Lq�O�gE�p�+�!�T����/WtGVѴ�,}����t��-���+�5�)�.�N�w��6��`,���iv?���=����WB	�y��~��<�ߖ/��c�Sy!�˻5������}MFg&��>��>��9�/��p���WF5��}ἰ��l�!���p��w�zزxE�섆�s�����ab�6?t��� �lL�5�R��(ά�����Nd4�hd@il[�)iX8�%e͠5\��b�yϞ<�,�Hb�&^�s1�g?�,�iO�"'9��i��6F4֋�̼4����g�s-�vW��y�q��[��Y#ʌ�Н��S�gE�|�i(O��9��Y�S�ao�yN�X()!F^�������
�����g�X$���o�f�i�e���46Kb��J�Y���U�H�D'�7��<!v��sY|_YRΓҞ��x{�V�?U�{�oT�_�Q���6�Jd:[o�f��vJ���iBl@2	BW��
�G�4R\R���h�e��M����=��QjL��Q7��|\VW�p����-tɬ�#0,»�P��pN�y��-�BM�Xr�m�>h�����K�%�1lUʵid=$י 銴���#������{	�p���3�J`�_d�C�B�A��T��q��p?*�e��c�0Wq�Y>��,8�[� Y�4�U��]�mdxyľ��Jl,"�4x�M[Tּ�53�e��ns���]�/qN1Ծ����F�*@A�}[_���f�Y�u������֜���)��6)e��رx�g$���8x7�/�v��~ɁSZ���(���k�w/�7�œ������Wr.&��PbI�_����B����9ҽ��,Ek	���6��6���!�P��Y�pS^8�=�DD�m�qL��omVO_��Xmr���"E���R@��ʶsxU־�A�N�:����p��ucc�۬�X�;AI����{������vu�y��a�t�c8m�Z-k��̮�>����	�V�	6cps	�?��"�g ֎9J��n]X�~���S�Ds�ޕ,1�I�!��+�����$t�Q{_���z�j�V�=�R�m�̚��V���4�x��к~��18�m��3-��>�RD';4�}�ToJބ!��*~ ��5�k��)b�P�7� i�dZ#sNnkm��5>�9+R���k���-��rb<�X�����*�XbL����9�!"�"v��#���x��r=7�Q�Y�	Ճ���*�}�����[*��t&j���^��Ð4"d�k��)���s�������b�	@d��Kd�>7+����R�\�?�ݸbL�����%R�W-�0� ���h�#��;È� ���H��]� (B5_�D�z�I�ю���΂�	Y(��cL����]A�cL�S�"�uh�b�/�)H�6V�m�����r��)~�!�!����M�"���Lk���L{x��0�Ԗ>8���&3�{���wv���r=��*�3�NME��¬zk��g@X�� _�v����O�p��nݙ�&����ǅ��rԬ��"-�|��>8����Ed̵a��wz�C�ݨ�R�P�$<���A0��gc�ٸ�ѥ���c�?[)��?F!�l\C������/�ӏ�^��ht-���o�r�<Na_¤���r0�E���6EjX�1kΘF�t����R`O��S�{�1�QR�i-~�c�Ƚ,Ƽ�0�[Y E�#�IE=SȺk��5��ok��1�^��0��_�
cPG��=�-�#<�	-�UM@�����lt�h6Jk/�X�����6�*��ב�Mkt�p�"׌c�!}���fMLI���<�:��a�����R��m�H<8`#٩<�p���1���ʧ�g�(Q�{��'��8F�&$2Q��g0Ą��yޡ����QTeY2���Z�C�1�ֻ����7�O'd���I����S�V��d�(�]i�y���;�Z|[�<�$H��x�F�ty,�&_w�HH��C{�����MnH,�r�-X�8��ɠ$l��4�NI�CD��Ex����Sg<��l*U|�ǡ�0���K�@�Pix^��D��om&aBΘ0����cX��T�C]��cp����**�X�E}�@>iF�@H��Vؖ�u�gpZ����ub�l��^��TtN�[�hP����;�y�⛯U�=�p�c���9�ݐ>�C��;��x�����c���R���#ˤ��l�j,a"���eJVPRRc�~Aqs�t�%MLN舄]��Q�a�)K�+��_�����]؍U��JY ��� �qSPɍ�	�`�IL�Px��\1����
	 ����ۖzj�N@t$�E�a��|}NР�k#B:�M�ڝu�?m��C[�K
�����tw1=��l�lǺ���
t��}ZÄ����N�x�Ѱe6���:}ٔ�:�������fȸ���_$fU��%(�ѯo$7��%Y�i@���'�Y��	�`ǔ���x��GP�z�،���.����&?��c�Ͽܴ�e��2���r\����0�\�Z�.|�Łu�XE<��/gA}l���4'x�Bv����٩�C�x��U�R����~��{�K(�k�8igV&f��9H�
�0mi9�S
��G��������9�v��OMA�wY��ȧ	����F]Z��@n���_��5�N�����B^��� �ќ�+b���ba��tc��}��}������m±զ�T<���
��jͺ������q<��f0���:�P���J��o�� 
�p��ʐ��a
Er4�OF�^�'��Z�-1�+�s���8��?D�3؀�ƾ"]�ˏ@e�������(ff�wt�e�������)W�-��0`�Z�Xw֬�}��hc$p���������h�JX�b������!&�ܔ34t��?��n��3߿5� �� ダ�]�R�:R��c$-��C-�<f2qef�3� �=�@J�j�`㐍����%qۗo�E�uk)b-&ct�1�"w�y�Ao-�,�6b1�"��i�D鿡��]���B���r9�;vT2@C��zω���[a�@sK�Tit��W�$v�����a�$_������t�����S�����~h�Z��׉>�?5kΐ~+�E��-��1v�gTKz�#�.���0�_��Y�h{$w�hෞ�~��<�!wg[yX��rS]���wf�uΞ�yi���k�-��b
c��%�qK�3�R�v�&"��d2������Ʃ����8�D�]��p�ѧ��-������>�B����R$EHKT%�<���u���N����P�%�[l�y��/c"���]�}�kc�3�I���;퇜���&0
�eƵm���r�(�e��9�VF`�V�i���`aE@j��b��;���z���R��m����\Ya�Gn��0�	MAzTT!u�&��qU��P)���9�B��И_�MC��l��
���r�6k�%%Q�!�	8�}#{����A�<������]�K:kv�$�ER&::Dt�:}������s0�a���+u�W��C�X=�}	��\�.>f��g����v����$#f�[zm�1\��7f�e�p�k��Y���e��y,r�g��D�-QsuE>��W���jAq��X*t"�uzW����*B�wb*� ��<Jʝe���B��/��Y�E��Z�P>:��KH���[�u��}��HH�{�9e|n��'p�~3��>�pZ�_��Fb����cT��*\Q5[�Ҝ|-U#��t-k�r\�,V�g���3 p���5�i�.)��t	������V�������Z���������!���(T
�"#MXx����Ӭ^�ޞQ��{�ك����@�mϛ��i"�Ԥ��I$�3�ڒ��lL�NH�c��/LxTJ=����~v=3w�	�j��}���84��¬%����LJ3��fQf�9]��;_hYf��{:�M>�).�z����|�@�F\f�V���'LH�=Qb(������Zf\��#>wx���rC�r�_X{�P���3L΁���T�����&�ى��Ͻ,�vQ@|�zGۜj��@04{7�E)[wx�� �x.����Q�p�a��f�%[��޸���0���p�d'���H��0S��q* �*3a�s:q�� zi1�!5����#s�հLi�.>��04�6>��ġO�`/r�gX�O$z�Y�����E�U9Z��RE��yvϕ��g���H�W��T�l�,��� |ԣl��
Q/ю��q����L
ز@qw���X`�V����(�D�M�{%g�{!�p��V�ݺ�4���mba{MZ`��;�'��V{=�w@{g"�(o̤)��H��6�VKh�'��9��5�W���ǳ�w�mј-��*N�N���q�H)��9(Ä��&����B\���D�g3?��/���^B�Q��* 8���2ĺ
��͊#�iy?��W�&�,�S:H����!���s8�Ɗ���I�	���ޤי܄�'O��ً�yc���U�������Kl�;��]Q+��ѡ�G�(��YU��͚��Y�kY	�i
��b�Km$�n��K&��V;`2I�ĲI�I�����egF� � Y���3�2i�wm3����83�V��#*���_��
Z��4��6Sj��}^;~XT{��a��<�m<����!q��Т�'�H!�yN{���W�z��tho
+����`T-g4{�)�3DVH�g�u�4�pA���%5-��) ���O��(��zV��J@�}�g\.f-KR-��4/���a�W�Z�X��&�i&ܖf���R+�
��T6�!8��ĤV�E7e�Tނ��s^��(|T� ���	�y �����̘�A�Bd[�ܯv���2'�,�u���((59g~������O?�@DXQ�̗5���#�����HN`���h$�b�|<hT�	��v����G�#Həv���9A��K-��t���=��]�_�>�G��o���1�\~��{XTL�9v�l�9�8����h�����\J�%�P��Q�j\-��	��<nLI�LI��'̲bH+G����+cF���@��آ�ϾYB�J�N�#�I�M����K>��� �c\C�x*$ �M{:&cd���������1�{G�#{�~ ��x,Ӿ9ńk܍��Q�J��ӟI�`�ĐrI4���}�A���(Kթ�Q$�ψ~�f�����n�z|���(����Ք�$�=9�!��7H�i��Iq>�"K��x���gC��U�L����{��Ue����ʍ���i���+�_]n�����GP֓)~��ӽ�7���c'6S���\�Q6�G�2�3��K+z�Vt��������po�}՘Z�u9�����]�;ީW@[�S���E�8P�Ù����	>�椞̏�ۀ�v�P0w�ݧ0�K��*a�r��n�r��$D޻��:N҃_u&�mH�V�V�%�p�~�3!�hn�̉��Рh	@�O��#L灁x���w��bE�?��a-���ElM�vj'|��nu�(�+L�s8��!��G�X7P�5��ފ�'������a ?���S����������Fc��)*I�u���m�r�sk�u�䰅�L���\|v�zHZt2���~ ��YT?Q���h^�HVFo��HCK0c����1�G#�h<}�[�79��˪��S���S3��+K��ʝ�9�B�#���=��$�~d�k���)��X����r�����֒Q~�!��:��8cJCKj�cǌݣku��{:��� �J-|D������'�Ũ|U�"����Y�G��o����ȷ�!A� ���՚C$�V�%W�7�;�K����{O�R����ɱ���������e�U	�Joxޮ�+j������:��a��?�����DA�"v�G�Ѕ!��W��L$Yoi�*�r��DH�^eV�M���Y�!�`S��C������6�$]J&�.+��ͪ�ET��I W_f3�mͰ-م~a]���?�Z�O5+�7�cbXļs���~`^>G�)�ݠ�\든(�V����~E�X���F��	�K�#�D��)ыiۈ���?��?��@��fdj ^�v�+]l�ˋ� ;;?փw�(¹��)�-�i.u�+D^��
&d�E����i���o�	39�ӧ,�MH�To�f�|Š�5�M�ưd�W�_!ڜ1��!�EF��%J���08�0��^�q��%%-j�rq{ Y��֥n���C�@?�2�h�F�T�o3D;����2�h9�{H�&�40�N���M�/��$���>��s��'_���t\���F����|ѵ�(��>�Wk;����}�ӛL��]`����d��We%�otS��կW���i�-�:;q�z�I�J���2�CҨ�Y�-i�X�e�М�^���b�X�u�\�j:1�Ȥ��<%� Z"� �6\�;a�s�8��Ӈly�(��XP����֘#��Z?L:��䑎�jn�;s���&l��� ejM�]Mj�)}"w��d��G8�["Bs��}CQ�(aT���m�r?�����$'
d�\^;�N�z�@�	*��DPo ���@W;.��R:(�<+��֜"������ΦA:R��Y��o�(do�+�Ł)Z�(iAX��Ǯc�
C��*��m�5�un1�G�t/0̋���Q
b�e�����C���	<9�^��5��;Ӱy<'1���ᷔ*-)��vn��`3�55G��n�l���$�����@q���du7a8&
X /�CU8{:����b!Y�JJ-��!�5�[��	����#�£����D�"bF����>�����̇�?j�K����{���MTN���U6���=)�h���Z�� ߜ��+G�L�@�^GH��n[O|mG��rQ(�vҜ����qw~7U��H�tn٫�"��ͩ_ia���$e�.pdʩ���àҬ�.4e݀��H�Mp	^Tbl-�B�-���+���!��[�1�I�n��,��J�a�F>��ꏬ7�[b���n�S���Xd�F�(S�L�[6W[�Y�B�\��[��Í">gK+��P�.̇Th��+rw�X�$���w�_� ac�#���l[N�!CG7���o����B�y#�ݯN�>�@���t�!�f�/-�	�Jb�"��*��Օ�E�B�0$;R�Z�Bf�L6ʪ�2ɺ��_
���Pp�wh����_����7°l�D>=Ϊy����?s��q�EϏ��f��Q�+�8�Te`��M�- �^v]�����w����T �7$�L��e˹ʶ� ���s�E5�0��8�1`)P�7*���˿��{�!�Jմ�I�9c�����,�W�j���mc5�������O��/��&�{FmE"�����&M�_z���Tע��w��O�N�OlY?ζ#�FJ?�{Yʲ!!_� q�g�SkE���#/n}-����u	8�o������ ��`r����3$��h3��4t�ȳ��\���߲bl���M>��H�VL!vD����S�.uD���4�}>Z;xp�ڠ��Q������A-�RJ�!����F/Y�]�҅<�U�L�?;���p���%�, :��z�\�mJ�G��Y�Y9���-�lP�˃���KخN��x�����Qo��t��2j�P�a��/G7bf�ܾ5 �5��T��[������\�r^�|����Yǋ�`�Y�XS����L���x�ŵ��Ngh=���=��{� 	�XO�0��riLw���a= ^�CT���������uD�S�_$/� �7�ɨ�A��J��8���2��0e�@HBX;�0�0Knb>�5|��gH�?��T�%!uL��o��Up���z��B�J&�>���y	SW9�_��':��Y�Z��s}Dn���b"13 ��d�g�Z��O�PL��r���uEw.��tm��V�E2q \.�Q���S�/��h��gX��9|�CqD+���gd�!�2JY=˂�M�ʱ#���=�1h�6�gDڼ;����m-�'��7ˡ(v̲,�)^���	�iDi�f�d�>H%.ţk�5�i坰�ud�b ˹�|��t!��M��(��nLեG����I�G�������8�
�F�S*��eh�v2A�C��|���sX����3 ��V�b�/k[�8X����W�S!�uCQ֒͟U����C�գ,%���.��i᫲�Q�~�(|���W�{�N�ݹuAG��Mr� "k�e�y���-�iS�w?��D�6gDc��S@��)n;1�j �H(x��~b��L^���Co/4��K���3�%[~⮁�U�;��k�~�7�>���ioBq��~����u�-i���0�s]��<$\n��#�ܥ4�-����5Q��0=��E��]3�:�Թ��Y<��A�U�R�EWG�o���#S�T%���!�I�_%z���ɰ��|ѰF�n	�Y�=A��d�Y>���^�hM=ڵ.OIHA��ܼ��o�?L�2q�mA�y�!�Y3L�mNx�5�sp �x�)9.���Ǜ�����k��A���IYBl���WeXJq&\�弲mL1�p�dP���M�j�ש��x��͆�l��ӹ���#�k{���=䎆K2�	��@��^�l��EPl$�2��c�1�<r�tJY�L���4LԚ�ޏ5��J!?:��Wc)��K�o2��S4�;�P��Gl�#��d��$��zہ����c���> �r�;E�LI�hd��$�^ ͛�'7{^�\e{��P�g���%ƀ�M��֚�;ϣ\9\됶��5I�Sl�M�:Ĕ��2�/�pr��<e�}������0�mHe�������J������"I����Q�/q"���&��NY��t�8���#���3����"|�݀�f��)�������&�U�m��[��\�Yƀ�Вa`L�~��bqO,�]��-; �`�<�M	/�hٶ��������0�A	���a� ��U1D��M�P-tQaS�r��sv�1�|���0�8�8�=�3a���k�	�wjdy�9�a�T���/��6ۂ�r S���VO~@�҈K���I���ѡ��μp�N�5���NQE��.��;����Gg/cr�E ��I�R6ư��zP>��� 0����(&�o��(��j�������I�N*pAh@s�,��J�	ǡN�F��ܣ�������� ���*�k��t]�`��zh�6Yp������j��ݏ�(i����bzߦ����1�s�Q�����@�['����?4,�T��s~��a�>o7{IFf3����չ.��VUP�a,c����yj̼d�n�~|L�j=�e������7h�!�љ�Y���J�&���>��)�<j
�D4�@�C^�ݤ�|�I�j��*B&�hX�g 2��"�)�"�,��G�ǜ�7N%���n��8�����cN��d�8qm��
�YpКO>~����D�Y����'R��N��쯛�ש��
a ������nLȉ�ֱ�ہ��ëD�T����T�WDp�J�"0�:)���,�+ڃf����S�(I�Ǵ�7i����DZK,*N�F��}�i	��uH�w��t�3�_z��G�����̼��U[:��x�`���f��(��B�\P@��R�dL�t�e�?\���ou��{�ϐK�; O�� ,WT���C]���5��+km�14үkL�C��5�6��Jtꉿ�-X~N�qAJ�K�.�\��%�H{-��~['�D�|b�I��,��x
ǆ��{�2t����A=x�A�A;��1�XXe �>��߬�}�dp(�9��۪��\ �k�S��������o��!���kЖ_TM�e��7ޡ)~�X��ǡT���5��f��w��Q�'n�0��-���UN�G#&E��m�F��,^�c6^�[�l��f�����uQ�P�@BX̎MY���O����y�� eA����+I�USY|B4v6�>Jb{`��'��<
:����;����{����5j[��Gac�X���"2K?��囝�_e��}X7r���,;�~��S�d� T�^_<��
8��b,cb�pR�1"s ¥�0o����y���⇹i�<���a��sc������6��iJ7�Z�q��*�E������@�Ԙ|W)N!]���9*������P��7���3X<��,;�C��<���
�*jM�Ⱥ!���Xy�4?I���	���g�Lj�tiƝ���897I�-Gdס�Ds��9��=I7�u��KdM4"�5��=��^�9bc�۝�^9��E��0��fq���[���k��p�����a�����'�H`I6�%y��F�P/�g���
 R�s��_���$�j���i��<i��,������q�?}�Ex���N��\n%;��k�r��M�����lMi	\�i���Í�ɾ;1S�d�̯����Z	�*��F���[os���"�ӂ.�����uy�����T��SBnct�u��!^��,�~܁+�+(�<��eN7��c �h����+$;��X���)��,�e�]�ö́�6N~8t!��b���(�D�b-���ڄ	ul�띈����s5���n ��*�C��x����M��-l��)���O5����;������S����IL�hf���(jw�D�W�)��Cƨ�#T1X/�zIVΗՍ��S��9��dx�_��O���EqZ�ؓ� �1f�=�~"n3���a�5���? P
]0���To=�������J�i�c���S�`�Pl�_�u�4�KrQG�v,�)���"0��]�,�ݗ��=�\��Я�)4V8�j�\1af3k}y�)Fъ���sFJ��"c��h��x�/-
�!�Ǭ��U_�	1��z,㈿��p�����ߞ���2Fdx������ֶY��y�7'H���X�)ʯ�U�S�l�i�H�pjZ����� e
�Y\��l	�j�8BaЩ�B3���
@�ŕ�΄�u����±oS�I���N�!?'B>dH.�GZ뙤O8 ��@�띡3T�X���v�1R�=�dk�.�'��a�J1}��x��u�}f��<#�]+*�p\I��&��,{|��%�����E&��jki�l�� ���'���"���wJ�$�w`-��{>����տ=a6&n�J�NS�i �a]P�+z�F/�)�	"�r�%ׯ��͂���L4������w�H%��"�E�BY#�«o9��*%�����r^g9�1���E��]��m��~�ȕ�H�h2䥧�(CS,�6�W��«�7�x^�� =�s�*jM� �� u��MoS�c�roC���zI��������"֐�.������k�����)x2(�Zw�߇x��P����.A�ƇR@����1�9���~���{��6��5Y�X�$�=��nL�Aj*�e����m�.4K��\�mإG�"���m����r�5���@�N\��έP�5k��u��831�lŕۯ�g�w��t�=,���V^�ZO��s���\�����<S��\��A༅A"8,C-"ħ��ul�A&٥_n�oŁ޷/]�s�ce}ЛV'���aյ���v!�40Q�Ē�(�_����x�Z�i�[�ZY8�J1rBDwG휠*�����N4Ҵ��w14h��үʮ`ԯ7P_y �Ѻ���"On�G�_���	���7qSA*ǁ�s��׈4!�����
�?��Jo
FPߝQ	 eV׮��o�|���u���8�YSI>.B�����4B�kq���g�a���[���r"�Qoѥ�M1P����ֵ;ի�wrt8鐞��<<��G>�*�%�svx�9W��jۿÐx���J�_�&F���n��K��kFy#K��eѸ�I��|����K�0,�Cý��O��ϙ�D����r��+X��>���^�SE�&o �1������Ψ��=,b
	G=������*���A\C`��X��{x/Z�3�2�̢��6V���L��
������n6x�g���QK`��x���1Kd�	I�Yk�|�b�M�s�����[p���h&@X�t�Y��W2�H#�������փ��xϊ,KHm�D�n�,��MW�/�۶��}A�5��0�*��O/_�<�C!����u���dW�V��Y�]^w`(���.&$�%�I��@�
���I]����EU�z+U�wTI?���*�",k;�����A����� �5��~6�-�;��3�v%p�'+l�2��Xʚ�&(�E�x�=���3pAu9�Ə;�Gq��_#0���^��}#�Z>��ÐhY a�Yh��J}�{4���xZ.�t[͹���\E;����Tv�y#����	Ѯ��8��0u�"��W�����>�Hl~�U�E~I)��D����OK�~��}������_qؙ7� pV��W^RIr0hÿ��Z�S�3{F9�z�YҷX�X�� M��`��>���M��^�(�\�s��o4['l��v���tR��P�� ���<ۜ���n��,}qՠ�=t�G"C^��R'��F��ڥE�M�O��הwO%6����{�q���Y�>�?�j��ØWtkTNr��_q��j�M��{xG;�f�{ g����bC���]�5G�Ƚ����:ջ�'��<��D����	��t^�5�T�W�e�
�'����+�Em��u�y�@ӈ��PV�q���YL�6�,A�*��|�0{��yOBE-M�w'$�Da�atS��!���VKX�g�G������Kȷ��{�|��"CQ�����nCi^R�Zr8��@��T\R|��v,cu���L��C�xF&�s��:�2R�Я��#L��O_���7Jѷtbm�p�*�w7F����%��d�� ;�p��+nb�?��ynoj�q�F�B��C�y]n�/	4B�.GQ5͗���y���fI��]^ Cّv6��6aa0 ��HTzo����5��3��lY��%m�u�T��k���ea�!�r:�����N,�q�)�a�U�#詢J�Úz��⠻0Oj"���$Ia�ve���O�}��E�*��/��5̚e��VA������ZmS���9�VJS�@��o(η%���F8���ֆ�Dʂ	V��B�}Ҍ׾��e1��?�"|R����+Oۗ�1j8z)��٭%�y�{��O�o3;�`6��<���'���u��m��0��Wc�q^F�D⿅�!�`�;��1
J=�ks��l[�lS������K
�V����UZ�tws�/ݯ��'������j0|��X��{��ᚄ�Y���	W�z��Ú\���Wq�i�m��N����g��wL(�ѠQ%K�Ɩ�H��v�dXM�R��i���
N��Ln��َ�ee���Q85�dT� �tn�_3��O*������p�a����L�/��)���+��J�Ν,ƠY�SP���L��P"�2R������e�.,�(7�����3�C�,ܪ1T�>UpZ/�G��K�+O'ģ��ba�;<l`]�赡�3�}�g����(nL���p���҈Xʮ�?�nm����>�Hk���'f������UYVB�_���0��$��0����p�=�-�UB?K/��:��O�(�*;[�$DX�G����fI��֎��/9ƱkY��N� +��>�q��/3o��[Z�6��V]��vg����_k�wY"�oU7�z��҇��[�#c����(k(v�����E�]QB�Yk���Ɣ=�i�EҚqkp��w�o�L�-$�o�J���pc�Ld��z">�N5�'0Z <����9l���N�UrX��5I��2f ��b�~����6���>#��ۯ���0BT��H �)�c�CF"�=�����=Cg�k�� �UZ6�f�TNª6T)�Xq:�ah&�¾��µ�8y��	�%Oe+�ҊY����9�A�bC;'�U�Y~/���q�0n���5�3��ʛ�6�n�=@�u�����8pi���9�c�p͒��ۃ�c�+Hޓg�p���1]�Z��U�8����u�.3.�1��đ��8g��bj�P�)o������g�=�w�O��1�TJ]��@Ok����Ώ:'��2
�EW6/˰!�l^>�o$��AǍ�*j�L�_@
�A}~�'Qq�����d���'�P�G����Oע����A�zCr?>��vD�8������g� KT}��j�WTB���gW1�e�XSx���<�`b���~D`��ܽ�KG�	�Z��+��¹�@�ņT�2נ�(�p66�s���=E/���(5��̥?v2g5C|�k�3)(3�]e�(̞����,��d��y�&��a�U���]o&ͮ�w�3��&5?|��;�V�O(<?w�'����w�r��D�	�ם�`_�		����4�%��Ag	��vw��L<��ȷ%'������wQ�@��R����h�Iy�Z�)��y��LE2��{s���U�E'a,ua��ϙ@IV4��,���8�u{`��1	��g��\;Ƽ�!����g��O���A�E� �B����|��e:�[�4�3��[b��I�Г�s(��O_3��H��1ʔ�����L�|�Z�|�^��J\�� 5]y��2RWN�d�x���~�&g�H�λ}f�즺��ߔ���*^������},���/W��o��JU~��\s?��P�Az��_�^w���t�Y�P�_�q�;$��P�\�Y�Nc�������N�X }�������"fiv_g���[��������N2�x�����e/��bȓ��9w�{�S�Wm��}�x��l�C���8A��u%KA���gwy�Լ�w����'�U��,��� �ӌ���U����cM�V��WK�9|�_Zt��㿳E�F���NR"p���F9�ʊ��Sk�8�Ҭ-�+��}��=�"yu��$�/��,��r��.��rK���	�?7fD
�`�`�^jC�@�;U?�P��T����yB��<��w:��I���aʠ>� ��&��b2qF	��P�$���|_�x���$\������-�P�~��Y�MH�-�Z>���%MOp��MS���#���Q2f����e]�i�o��[���B]Ӯ��/��˷�����t��v]�E��(_q��k���̚���t�`%��+#P�.Pg!L��
m�Pr����"�*������i�Y�:�Z��cUsV�J���)`�b��j(���Mۡ���p�c�8+坨P.&��:�zj\n|���N��X���}����dϡ�d����e,p�k%
jᇴ��|�6��G�z"S��C1/P�E�����.�4���ԓl�p`a��e�[�A.y�*Ќ���o!��o��w�b�;��ja�����.����%���	к�g���
61H������n�����~U�+��A���";z�;9c�{=I��l�O��pH�i4*�3�*����6l/���V�������Mv�J���Dc��M3Gi��f��x{��S�ht,��>v��&�SX�I�Ut*yG���,��!N�H�o�W�:�5�e(��q�T����@��|��B��P�y�-y��wHrK�[.����{  ���É`��:���2B��H��v�~��ٰ>�_j�$��CLQ#��衿1���E�\�J����`�,ˀE+>�L��k�����/�u�����H�F��iGo�Ѩ2M�򯖆{�Wk`��Ag軲Pt/-l����fLa��od�ek��y;�6
y�-�.�0�	M�#�N�Pm�K��k���Fp 6X�oY����/��+w���_KM��/�� |~�4�ώ|�I�ȉI�4J����R�y�F�����H����^����B֛F�9����d�\�@��7��68�),�	xd�>3���iK��]�[-fws�&����$�7���uզ������ż-�3h�{�}(��K�e��i��L�� � �;A`5Td*�i�<�fR�Y�/�����p[���9i�+�:C��3�2ј���mnF�D���&�����f�O�0w&�;�_���I��3�a`�}~�_�/�՗�\ZO�]���_���Q�r���Ȱ8���kT�a���q��jq��á4ph�$;�8�\��W�(d���g�|���^��F"N���Ȇp�*~�%�I$�f����7�nt��S@��8T/�.�v�����[�K���!�'͙���=�}Ey߰Z���}����s;�B��ʢџ��b	_�-݉T���+��ϱsB�4g��3�,���a2���K1yBn�Sj��J�������!`l�)A��3{���I�0���}�$�C�j���S��p��8/����VX�A�Re�$Fu0�U6+�*Aq����CR�+33>�i��/4[�q�_Y�����g�&�[k-}��w¥W[��]�6�*n|����Sҙ���u7$�k3Iʳ�|�	Gd���kK&�HN���@,/����͗猂|��x��&�B�0*��n7�o5vJ�k��
�P~��Y�7��ހ:�����)�N�p̝;���ގHd��'�i9�Wܝ;��^-X���
�P�+�<<Ĩ=�?cMɻ�8�j�tX٧�{�1���p��.C�q�Z�(�R��9�cN)
�U.Ќ��J-�`�����ڂ	0T�Eh��2��z_�#����\�.�p�3-��G��)�%��<���c��;0<��] QU�<��U[>�泚�+�HܤR�7VpOxy9�k�π�Z
gDj��6�i�ƅhZ�U5��L��&m���Ld��1�o�Y�Y��)E�!�%���* 4�oUc)N��<lc-�����;+�G����;���!M!�L�%!�f?.<Y9fW���jL�toKHԦ�n�2Sc|	^�Й�u{�x ~$&�~�RB�fEg
62������ͥ��ƒ >�Il�l=K�1���3F���	�3h��@��3�̘-A([�E+�v0�=,��`g�P��M��r���d���L��
�ͤ'���"�mT��a�������~�7�
ӣ���Ȍ1�֪ @�
4B�Wd�{��@�of�e�IX��7;3�m����Y�m�*��@��}hXU�_,��K0�� o[�� ���@���R/f���h���2�j�터��')��/���3n8�#�?�By�m�f��@8���	k�q>�&lƇ����l3e��F u���s��N%�?�#-��<8��Q��f����J���l�Q�.�s��!q���%�
���2��l���G������B)�<�Q��-�D�iiv�0�O�3d6|Wr���� (�����p�2�)a��D��B�>Ж�L�T�S��/�*�ro��û/]��Y_\�M|PRV]��	 �'����oj�ls���[j�jDa�Z,%�a�Ha�a▗�xX�6.�Oz��qW@��)g�R'�qF>s]^&[���7p�^��.Lb)�t���8�B��҆Ry�K��$K��G�+��ׯQtɓ8�i+���֣���SW�d~��3*I`���d?������Ӆ<ҳ%3����$�z&��)����]�ϗ]�I[�[�o�N,]��y��$��/�7�����RO��VDŐ�}�o�F�����G4O���ή@\��4�.�+�X*_|���ۼj(+>J��� �T�~��������?��e�Y<Z#���,�j���]�G^d�򛭇��c��5�^����>��;rm����'i��=nZ%�!�S�)�x����K�`x��m��tUf����~`�oB��{��ҕW�`�8����d����#��i�[Zc!��;�)Mé;Z� >p?�P�(��Eo�����v�� x����bn�9>l��o=�xоN��~��«�n�3�+�M��
�?�����L ���l��/Up7��O�ݵ�C��|��E�]��ߟ9:�[��f]T8��������C��x�2��D���A�9���7��L����A�Mp�P����M�k��]B�B#���������w�Y-6�p"Kv=x1�QI���
�.S�����kR]!r�7D�EVN��ֲ%��P�˳0B}�?΂M��P
�"C�i6������{��)�T��s�X&�O�K,��4��|�~0���Llf�ʗ���[?�g���]�:1��G-1]���H��y�o�����H�
��۟g=�V$�Hևh/�wB����[��İ���4Uj����3d���L��ݘ�3K�@�ܳ՗���tF+�W��~��S�� ^���tM�<j�]%l0~۝��El^ �� Vu�Ъ��$A�����K�����YV��>�fO�N�:��U�Miy-ӟ�-ٰ�)؊� h:�������rf&z�=D��{ U���������d�$I����{.��{�R"ޝ,��@ז8P�G���P�h\T�,2�͸,[��X����f���l���d���{�ߙ�(\��c�2p~ e��8�$|[x��s��7����	
�D���rn
/�����b��*�^ǽ�}��<f� ����~�
x��ф�Vf^C[�ݱ���zhro�5Z���X�J��!;��[IڽA鍄�4|P6C!rHF{˗�?����CTBg���y�ry�J����1z"���wܣkh��םxnÒN�������i/D�O^3�q3[-��'�{Mh� 5b��Jg�<��\���Y��tr������r��^�WeAr�	 �	}o��L������l���_�ǀ��6oi�+}8��`)Fա3��׵�=�Qߟw/�Oz�l%�v�$fA�U��q���6��TT�6,�^Q�ຐ��zeP�E޿� ��1<Ý8�z
B�@�#���}�8mS� �(��@�%�oV1�K[͵'�G���*�n�!�l����$�tG�Q�)��Zr�]�h�+Oy�=nWȸ��v��4I��3���{���/�	���F�c9��0�m�BD���Mô�	<��5L�=|���@�o�#�(��/C<��o�u5�5����k&�~j]�k���uY=Wta<*��A;��xhiM%�a���\�LL�������*'³	�Q�[{J���9B�{F�^���$�o%�{�����p�G䩥DTXm��d��髳~�,� P�5T����G�u4�Ɨ1��Ǚ�=����/NˢjA���n�ь��3IRg�S~a���p%ķ[��J�.����0`��Y!Yz�7s�1��D�����v)Խ��#��\�Ș��W'[��~}�Q+��I�a���Z�p�r��l�!@) ��^k��~�ű�<ou�K�E/瀰Yl]�n�7���=��c��-�i�Qe�Nڶ��W{�t$��&-�����s��Wј-H�������P��+єR��_�W	G�C�1�����|�סЀĆW��{��;�!E<�*ol�_�Ly�%�`���<R��眈��`�2M�`PI�2F� B��~FP�1��%-��V�����.�*����<C�Av��
���ǡ��ՑJ�0���&�T�z>��F�ɝI]©_(�o,Y�b�zñ;���.	o-��+�HXDg_8N�V���Y$�TM��T1��B���'¤��u��C���'��"�"�[���i��0�ş!���-�%��j��4kSa�X�S�䉌6�8"C'�	Z��qN�L�Y��+�r��U6�V���J(��_��Z0&�e�]�r;j��`J6�udAܻh�?��R�����a���߾/8RNA��	=bڿU`�ދE�\b5�����))��L����{�=����~ad'�-�U��.1`�3u��;�#Ϛ�����&���}�[V?�\�pѪ�#N�G_�MT��mG.dM'�t��MtuXQ�������BbJp������5�̈́�3���ж@����V��9Q$M1FU�L9/Q{�����n�����M����؆�C�0����`�GOB�\B#���4�+���H@���64����f�D�b�-�!&ы���XhG�BeCo��]:3���I�Ye�G���69��k��D�쩖�[�Ŭ<|R���	
f�h����O������(����j8�8�"�f�C_�c���:����f���������h�&��TP���X�~�z1f𨓸���Z��t��Ȝ�0�����z�8 )h�xJ�h}5�y���N��ƿ�iO�^u2��&��(7e0���K1�	��&f @q���&T�;�e�>���Mh�"i��:�605a��_ZWr�,K������|dP�rXEC�NVU �v�O��'����C��P%�'M�ۂj6��`7j#8�C<v�B
��@����^y�`p��8��y"�Q�r�1_eB-ʑ���)5�ؘ��5}~�)N8jK��t��5�^�Uzk�kGd[�a[)`'���=b;���	�c�;�~�� ��g�/4}9L�N ���P�<�6LvˤP^h��ߙ�,�Ẍ�y#9VeQ�E�yt�ּ�F��q7wC���2m�)��� ޥC�L�h�e����ı�ʓ��R�|n���<Ѡl���l�H��U�c�Ҷl̎.ڟZ�jz�;Gq��AcX������Ģ��g�2��:,	�6�U=��Jf���!ٹ��Vh�j؜���%�;յ']�m