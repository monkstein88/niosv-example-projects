��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a���V�h�x�Y�x\غ�;���rZ��H�Z� ��]]k�\%�^��|���_4����欌-�}:kc
�V��p��"��#�4N��wx�t���8k녬j\����cP�+�~�V��mGO��������*�h�B&����m�$��+nuUv�]\	}�G/2Zɟ� q6Fe��h!Ǖ����R���vK��]��Yd�.q�o����r��Ɏyǔ�����96$٭��M^���ig�P'/���+� �}5����E��[�"� &�����6]��,�?F�#���٤ܨ����?�t�#��V�hQ�}.�2p��|1��^^��|���M�����\=��+��;=JW���F�my@lޤ��z����I;*s;v5�)�E.ixR�JV5CU ��Ȓ�Kd�W�4��n�1d�2��?����s�N�]9N;<������d)��Ć���s��QE�L�;��
z�j��`/W��G�4�W�����MB�zR��<�Y�k��A~�|��׃^~�&�/j.�z�^J�Y��H���z�D��2:B���]����SLT��Y�e��bM7*ߍ�!O��-��,�^��$�	 aj�1�p(���fb�\�\�����"=)rA�N ���ࣾ�Qw�Jb�7������}�j=����f�;[__m&u �ˆ��nK�K��hu~��3���7�
��ƫ}���Q�3��f��ʣ
2�F��c�f���0jB��,P�}K�3�ޔs��!��$]q�֬:�oy������zsO�z�(�X��I_�F.�sT]�"��K�����v�����C�w�ס���|�M���M�w�z�z������tl3�ֻ��q@���K�����W:�jE�lf�H�X�_�2�N�(V�}�F ��\jI�ֱ_R.ѯ#�����~��;� �H��[$	k�C_rw>�j<�(�57�3,�L��
��M���~�V��u�*��)�N<�."���3p�I�fE�h��6�B����o�
-�0��5E�E˖`���s��a�n�z	(���,�	ȥ�ð_�t�����g`8�c{B�	s)̧K$��t\��p���Knj�AWAq�����O��]���׾�
̢�Hc�V�D�]��E,��EJ��K_;w!��/��v3sp�Ot�6�M�J�E
����z�#��k���o��O���dP���
|	]�2�/��?��l�������������x�P��-ǥifc𚎹���(#e�@Ih�I�N��P?&H>>�w���0C0877\Z����S����+M?:��V(���!�>[�0�)�]cnl�|�"݄�P��ԁy��bysϨuC@|�`_���`�钸��n4<ߌ`}x�:�k�؍x��#�l��ck���V���:��(��,�t�5�Sz�#�YK=P��K��*_)xfeɾ)��rR$fT�	��.��ʡ ,����� �JQ����~/�,Mb�Zdv�J_ƘS�w�����J >f�lm�=���	��Nc@Ο1;n�	��v�{ړ��;3c'��٣�����U����Z*��;2�[�x��u�����K�����(-O#bR`8Pp��O�����}��³���}��[�:͡��<ߋ�[l��$�j`o?jgK�v�  �~���A+ؙ�����-0���>�@%Ʋ$9ؖ�8c���L]�}&j@>������0�0����P:�L2���R�*���f���#�~	���o�Gc.Wi������LA<�'	�A�z������AH:��絞J`���$��?��dh�8gm ���*�
�Զ�����F���T`�x��[\��]� 1c��@������o�Uk Q�����{�y��&Bkuj������(H�UU?�)��8xכ�:kե(�����L��Vl'�'��%G��M�VC�z�:��-��Po�k�[��TƘ찼"]'����c��,-,N\�F�u������w`��!�sGB� ���heoHp�q�Ԛ������]f��5�]�O����s�պkU��kj����7&�c-����'�R%�lBp���;��r��!~�P��S����'��L�M�4��W��y�ʄ,�B�5s͍���&�9�X��ڮ4Q�l��x�@>�
��_�~j���e���K�q����g���o�j�C�� ����L(s�]0Q�?��J�BB<>�lM�dRlE{=��A�S1to��}��=������c��%��9֟J	�s�i)����C����<�`ͨwí����|���r���g����q��jPK�#�]��? �^=p���=�@�����Q��b��&��J����3�v<�I�H����yX�eS��P��� ȝ2_�냢������QE�;�7J��ڤ����_*W�R^N{�<}����&RA�=����_ ����(�~��K�\���R�M��O	;JK�Ż:H�/�P$���%f�o�V�~k O�R�['��}��e!����1�j�RˢN�p�7��C�^t�P��RL��dz0��YG�޶K�����t1v���������y$_;}]cE��E�8�X1��j?��B;߄�S��&#�\w�X�,��ZR�ya��y�ʭ��4oq �lo������}�q�s�c�*P����(���$]n��u)����7�Ҫ�����rh$a�Ka����@-~���&�߁TON�Mڹ �e��x�0C��wF�Ջ��\iB˃�b#���/I��/	�8�ۻ��d,���:
��zPdEſ���7��R�C<r_X���q��}EуMx�Jȇ0�:��	5플��#`������S?� u�����Sr����$��OPz��M6��~��S<��@|�@��T���W3#�rl��k ߠh�S̘�
���i^]0�lK��h���Ҙ~�B.�<���-��%� q?�5JO�i����kAM%��h`�s�px��C��l�j���C�F�*���5�{�V�ho9z^�6W[Ը�1��Qm�Y<!�&�*����CC�	C�i�z�a�J���ٺ׏��S�W!��Z�墧�L}���Qͽ7sy��]� Ǖ�,BC��,�[F>���Z�z|'2NI�Ё�>fk4��'��*9����L�v�:r��Ӧ�����x��L��HFG �	��\f���`�H� n�~����577i�*v�#���Y;�F��Mv�>����-�>�%��^���,E5�j+��Y�h�No�(��F��y���MUǆ�c]��$잍}��|]�sٖ+[������\c���	A� ���:�h0��	͈量����}�C��N`2B �pV�uV�Z�w����j5V�S��I�N
D���$i|��Xe�Y�I�B`�>��LnA�x�Ϛ�Q �:G���+�X�S���%..w#<C:���(�]
L��w��Ť`�����MHrv����J-���OL;�&pm�����8�&����{z����! �B�G
�l/=pI���@*"��g;}��0��;{"±mU�=�V�6Y�uJI��J��]/t�Q�	���!3��7�8�������m����4ѻoM(yV�����JzH���I���i���n9�S�ၚ�������)E��?��7������^�%�Ѷ�o ����e�L�ڪ4-0��q�
�}�UMf��`��ۧ3�$w'�i[zl��96����t��[�ے+��I�@Y��OCc=�ˋ?7�k<����|.݇��x�4?u��0�_!K�[��t�YDk��.��P+"�s���3}��І,]��V���FĦ�RN��N:)�����S6	��JN�| Xm��p��e~��X�����I����V#+S�<#�e��.o��Eд��iZ�KD*��tocǏ`k�����ڧ�I���o��$U��(�,�T0`�{���ҙ�� �l�&�j,���kGv�sf$��f)ZǛ�''�x����Oc�8i�	�G%F8;̈́�̪���BI:{jzR�S4��U�g���]u�E�P� ^�6�2),�� I�PU�T�67�bY���ËC�o��