��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a�����{������#��j��{��	?+�g��-��"XSʌb������;�b���/��.v���9�C���g�A0
��}����P((ޏ�Ő�����d��T�f� ��?>�ݿH��L֒6�8��.�~g��k�B+���ę)<���)f�~�7���
Bπbv�-ˆj#���`���sG���k���O�'3���I-��D�ʉbٰK{L��^�D#-5���#S�1���" �ã0� �[�~�^T "{�(�<auL�%�02�#~3ޭ��rsm^������.BR�q���n�G?�r5�?�.��?����+�7Y�l�?�� ��(f���p�Ĝ'Ydq0!W�G�e���x��.���|�t�>�⛇P��6��<}�2)�����MW#�G�˛S��Y~oK�����Cz75�n���U��Z���.{�p���WL+ѷ7F�¤q�w0��0{�����off��~4�����.	�/�Kx&�۬�����>��O�Mi����F��3OM���A4-<��E};�$���m�<�:WA�g�9NԦ��g�����ꎮiֻ��y���Cm�Ct$� �}���*��`]x����죘�h�b�;1n��������y_�mO�y\���f�z���M�C<��>S�W�ɗ�@r���T���a³L)f�i[σ�t��A��J9�p{��	Z�S�;S�=;LD��'Au-z�-�˫!�x-�n w}��Q��ʧ֔��I9�C{7�]���BԀxlBV���S��UEv���R%�$B�|h^��h�WsşĀ�9����J��߶�<��M�����#ᭋ�11�l� �U��!2�f
p�t��nit�6�?,����PYF8�_q��ާ�]�W��Cv��$��I
dk�ư�ov��e����{UUl���,��e�U�{��Κ+ز��8XQ�*w� �v�>�X8��5�#8��_|��A��=�װw��I��b�'�bv
s�hײ��+6��9�ME�4����Y�w�~���\�	�W�%u
�ś�ҝx�k�����)��Y�м��l�:��'Q���r'��t��&�jp�7>�=�/�\E�xbg#��,d���0��������p@C��v��Q���gɍ3�.�Q*�8݁zKG(6�����#��A���o�	$�N��n��0�C�lb}�s�^��hx���[�������'+F!�#yf���c�tPħ��第� q�� 㫝'���}�#�w�3"����!U��_�ز	t>\�+A}���P5��0i^��8_k)0�g��ώ�"ʏb�ωUh��v��6�7I��2����t�H?i�j�Y��J�*�7�p�����Hh�D`������6n:���Q�>�#���byז_Ѓb�@M���$���8_�I����X�;U��E/�5XZ��_
UH���vx
�@.��Q,�_����P(�_�v��ר¼�'8(��OՄ��w;OOIG�8�&�����ފc�)��k����]�X�����j����]3�c�U��`=qޮ��C���(~U��r8�aU�v�$��a4$�No2�S��lҭq���E��x�ӮC-
P)�X;��P�e袊rY�0��9��C���)v���4����.�3̥[���E.�Ʉf7�0�z�@�70���Ǚ�*+�T�ګ�v������;A3���X�c�$��u�a`��$��nDG[N���o/;J�%'��B8+uX�L
�hGk��M�e9�I֖Z���YP�W@�b�����_����U���f*;;�5`J�II�/X��:Y�q��W�x�́r�.F��+ln^�3�M�XQ�Jw�16��Xǲ�-4iiv��������ޅ��G�3|�ތYǘڕ����b�h�!�:�ҷNM����2!�1�ZS:Y�n��i�����u6�VZu$dV0����=���������B8�{x�-�M.�!�,+$_���-�g1����7�IB'u�F<8�dG�9��O�[ԂF�ֲ]�K���6T� k8؊�2��H˪�y� ZJ�d=8L6�]2�{���E��\~���cI���SdٲOÄfT�T��[��?ʭ-�N��[���Xך��vt�H�/�6�%�r�@t/-����]$WF���E�@3��zx��δ&&�T��K��!������)���.ꘔx&�m�tG��]�I���N��p~�-B$��рû��I��Mg��Xdj�F<�1E�U~����rnԚ�|�̗�Oޠ`�m�y�8x�s�4�;��u>�f���c�b�!�a_"���A���6��$j��muǍ7�)]��ؗ��\��7yC��%$D~\B���s���g-ޔث�������l�G�+��q�UK�ܠ3R8��"s�U7��sҗ&��.����ȓ*]uK�v;����D��������:g�؎�`Fh㻦o����������	]��"��YR���q���SܥC4Ż^��?[��)�ߌYyj>[�43A���r%jKAA*�F��S*��n&�(���$z-�g��GVzRHr^��i�}bC�y�y#\�����L���<�#x����˔m���f_��w�9��o-}��ɳ�6�,��H.���AO5�������A�;�@�������mSd���_
�tp�윽ٯR����,�L�������hv��mee������z�ǰ�Kz�G��y��ˎ�rP��Ht0OƹM�Ң��R�h�$F�d/���rG�A�@#�Goʟ�!��KR����*U���;�u>y:)��� ����e���=w�=�[ ���tg/��g�B:t��gi�ʂ����W�Ӑ.{-:n�I��fە�b��O��R�As�"�H��:�>X���"���Y�u�]���\r�m�p�qJ��C+o
Np+��|!#8���H2�"����;���PR&�W�_�݌zWޡ$��S]��8C�m�e%�/�LF-/����,������Yb]�3V�Gk}�)at��ȷ^�t� 	�e�p��N���k��l��n�=m�^	�1X@�)�~نj�b�`�R��/@|��Yk���|��^YY��8ϊƕ�%}���"[�и��$��ҽ�2��G�xr��L��s�⿹q����B����L���e��R���T$4�"���0�o�s`�]��,������~4��:���L8@�����o�J�6Rtұ��>�0��N:?�0(��-����[�,��X��8e3�6����w���}�M�[�#"Yk�����)?�'v(@���(8�)j���^�>6DHYs؉���r\T������M�5'�&p��#!.vMk��⣙�{t�b�:���òČ:'?�sC;Y0��y�iw��1�w�F������#��C"�8�7��z~�>�?�cv˰ݸk�*�.U���VKUljw��E�}#�Rs�a��	�rHl���=e2����[6_�}#�`T����#���i� �2'l?D�Y�5��3���k�++bn���A���Gz���`w�����&W?HE}���L������Q�AA��}Y�lDo�������AU'�,v�<�e?���!�U��0H��s�X�UE/7"� 4R��gŲi8vx��Zt����~M�����������n��US���3^��w�Z8�mW�-A��l��k�b����_�Y/
�-VG�u$�r�6K�֛`��KEL�s(~� ��cR�2�N�H�����Yf�#<�}rIs�~#�A北L���S���V�X�RggH�!�y���r"�4�Z�v���L�*�wQ��u�A�vѩP�&�h�`�+�ʅ,~�Ω��Պß.�c�3-)Z�O6�qʓ��"Zbv�S؅�<W[���z���)��ouFoǣ�y`����]c�M���.���(!uߐ��E_�$]w��Rϗ;�AG��A�~%��	_q��o�U���>9za�)��#�G���!,R��|��i6�� ���x�sYgY�J���w!�}�!��o�*��[�����\``_K��3^$<�E��x�վ���,	�@&-/	��\ �xMÓ(>֑3�;(�C��U��G0��x��;ٿ���y�R��ES�Bt>;�l����<�l���^�u8P�K��e�A�!��<��;���+1�<������A��8u�$~��lJ��ܺb@7���K�KU�QL�,�g+3�Y��z��I9��h�k�Z���Wt0����]��xa���;��DΪ���k5Q\�73:����8Q������~\���Ϊ5�	�AD�]E�b�i| �Յ����j3G ��\�Jrh�4�HL�Tc�O��0½	�a�����ͫ��M��6�mTG��A��ib��M0�컨sm|�z�b�[½��>#���R�����c�<~����`ѷ�A��`�
�B�x�8��Km![�۠#
X>��P,�3��%�hGwu�d̚����7?���j�ptY׵�����V���5k��L�q'IC����=R�/�9�I��"�}Y�WG=��.���Vb���JF>�<�Mea��P���� :��]���W���죯����G���Q�8�ϻ*�%�a��h�/�ߠ���Ρu�/<�%cEq�Ŋ� !�<�z�B�ʣ�m	�ܘ�n�k�z�ocș�o7~$���k��:T? "�.��߷&wz��Yr��f[j��+���g�v����Ms*J0�PX|/�fM �7Y$,�8~@do.�od����,� b�{�Z�h�������-�ea4�GXIR�9��Bˣz���])��9��~�l���oF���+��݁j���>gek���ґ[4���j�	1j}~���s"����$�m*XJ�h	Og�h�
G�<�/I��t��B.���_����
�*Sb��K����b���W��9�{��r��?��Y�W��W�x���|�P�g��C��T}9|FD6d6�\^����N�S��c��/p���%o�u�ۨA4p�yBc醘џ��=�����3���6�ƹ� �[�ʭ��m�L�Fv�����&���!�����fK��{.� ����L_m�^(@`^�1������x�Rҥ���,�#��"LHȵ́.g{�ֲ	�I�^��~���/k0`&ˆgPpwڒ�F�*n�I80husְ�y��*z@cl�8+x<��xl<�k�ҥ�g �����9˨AД��3����&\8Dy��eb�w�-��]:qf-ʗ�ֵ���q9S���'�.m��>��K�Y8�'_d6��QL��c4ܕ�&E��'L	^[���R��uAwrTPǏ����e���P7��e��Y���߫c����gA�$Ɂ.�B�W`��B��:jXNzBj��M�2#��1�)� �huբ<�C�(բJ��� F������Ի�[��9PQ-ҐLJ��jp�#fGT�3u�7wcnr4Q5*ͲQ׳��6�m��h���6z��&�OQ�@�S#�2��8�A�#PU��o�ƹ�q�٣2��$A|{���h�+��J�6Nc	|4��0ɾ�OԳ ���!�邓/K2X�w��Mv�e���a��b�s��\�rXҽ!�T_�a��F�]\߸�S��"Ga�(��Y�٦ �<�$W�����hEc�,
j��K&�Āשv�L�0��x͛�������ع��3 ���L��횾���
�|��\��^��]$/蕹e���g3)|��W��Y|�3�h�NF9�f�<l>?Y~4�zྃv�.[������.�f�V-�,>���|֌��X�U�"��C���B�+��>Z���U��-�ֻ�I�0�p�li�+| >�?lW���<*��2{ڴ@E%[	j�ڼV�J(^�^H�2�G ���c��yJ�Փ�`�.�*&��o������� !Lm��,-�^��/�·*^?~�|��\w��t����s�3��#p�6��lX,���i��
�!=��Pϡ���0���qQ�T��pUej{U�z��scC�R�I���Sfsp����L�ڃ�E��v����_��d`���f��'t#Bgnd�<s�]b6A�vio'��?��0w�W���\�t0�	ͥ���e�Pe����ɗ�
i��$����%̀/�RO�%����q0 �aG̕Õߣ�\zW�N\I-�������1wĪM觴�C�޹�Dqo�%%"<�0���O{kޱ�em�g�`�,3�vד$ū�!���GDG3�(s���B,]�$�)ͩ�_(֧�D�)E�s�nq"��Q�E0h��|e���N�N��n���1U��R�l�'3�ֈp����CX>d������h�Vx����~Z�l%(3 7	��~k~\d)U�P,�(�8���M	Ty;..�9�/����_���������!��G�G�U�x�����f���ws�6�"�3~��_L?��ɨ*�A\6G[�"ff�j�m,x�M�&�O���n��t�=%r���ъh������b*1x^Fx4P�t	�5�l�~���]дE���h��4o8�u!�%�yN)�wɢXJ�e����8�{�>������u�)��z$՞�	�K��z͉`RHَaM벧����]�XJ`��p�i�f�U��mַ\��e�'�]�:\S�t���Ժ�|/_ r�a��M��"|�FxT��Ҿ0O��`�kq*0�ւN��vB �������Kr���D���W��|Ir�d͝�IXS�Zǖ�8�8�
N�E<����5Ì���ɦS���T1VC�Z���E� ��ӕ����!i�.R
J���t2��{��>�y�I_ե<]��؝�X���i�3��6�t��%��^����
��,��r�/���ؘA�t����o�f�cp�����	I~�N��F�d	jh��?��D����_]H$ >����J�% Urv{��=4�r�p9��,1�+Y�K�M>n�湳-��<E-f���'}o��VN��c��-�C1���&�pb�&	��"��?L���A&�0��;�I�
�O�
��# �E��}��G����r1��F'�-�&�ҋ�Z���l�q~�j�`��k��=FI�cpU��~߼����`6�R�;Ɛ�����z�+^���X��Ä�Yp;�K՝P.,��p�!@�,I��=� F.�A�V���|�o �Q����+HsH�Ȍ��g�\��Բ��v������a�Hm-D��וkc�v��KmtDM�4I�RĿb��`��ͣ`��5�v�L~�u}�|UD&iހp�ŋ)Ϝ�Lz,c�95p���&�} �-kl����sQ��@��͸�6��hFT]_Q��R`>�+�&���6��O�"��ݖ���J=�c��~����۠Z�Ef�$��:���Z�
��]�&?���	��鹬��:5����JI����L5�Z��ާ*}^�H���_�Ax�	�����OI�\Jy�8��t�p2UG�N��,B����Y��c��w/�4@��u[1ơ}-�H�6�K�8eg��?yp+%5&�#�o0k�Rb%g:*"�ޑ��!�Œ��9���;k���֗���)�SJ�@�-�Tv��t�V���n�/�s--�p�Mee}�9����_|�#J�D�X���S����s-�	q��*^��a�������]�j
0�\ꑮﳣ�..�0��u�t�C��Ǚ�+%�Eś!��z5]�YjH�X��T���m�sv�z+��*����~�z���`vDR,����y#KcJ��V����p�y��eq�c�)��x
 �X��i�봥y.����$�hjO'�4�_��bSК9?�%���3�:���J��m.!f1������(aPG��z�\?{�Eơ��&Q@��ϐ�㳭�	�ɦ̽ڋ��9�e�]�5 _�:#2^�3��&�;��>88�g�z�g��"�#�X��+�.�0���۽� 8�t<�LP��c�
��D_vflDj��<���6x+�����v�
��D�L$�/܏K�gB�/dr:gpW����g<30t����~��x�K46}��~�U-��Bб�y&l��E|L�3N���R����,t>.DY���z����W���T��}�QV]e�:�����{�£�C>	��\W��ôB$��D�M5���)�V�& N|��ư��uK8G��'e�t&��o�L�@������,�#/��(���~Z�lA{ssL�*�I��n��qo|�H4B��=����G�GO*x��[��
���1#h��#�Z��������
�B@&"zſ�)���svͿ�����Y2�����}ADv�߰�+���4fbf^��+b�.5K�u�n�)C�	Y����&4�oޱ��8��?u�ĭA�S��բ%D�2�Lv
��ǧm�-�j�1Z.�* �-"��gV��)��4 ��:�%]�g�bG��������N�2,mz+	�����|<�6�
�w��V��d��u�'}����w.W8(�y���_�
E��r,Zjqԍtr�4Or{�F'3�g�Z=�
��Au�
��&{���.�\(:=q���T��1mF�Iv�P��f���ےY��=�a��)!}Op4jş,6� ��bX1����	�.��F��_�y�z�<�k	�ԉ%�]��j�ؤ��H��3)��B��S>)8����zujrm���]jBD�.�0�K�C�b_�ntI�so��8�.('}QP��%�}�
&[	�c�u&����?� ���o��wJ����9(� )�������}��'��잢���N���L��t��\�1�ӝ�1��cQ�N������.ѥ��w~��w/ֱ*z6S���Z����~I*���i�[�c�x�;���[n�>7S�^(���Q?Fq�K�HӺ� �w3�΄���2�0@;�����q4,f��o��0sWC*s �P*����N��&�"����v�"bqr�$��7!ǲ;��yLb��k��4�Jh�Hh��\h����3"P��Hn�M�~�i� h���,���,y.�5"H���Ø����x����hj�-����n1��Ƨ�RF۫?b��V�
EQ��_k֗@��r�QC�t#���i=��;�H�A��/#R��-&w���좔��4���4���%��s�kZH,_ȉ9�闓s���'tBh�����%����mnL�p%&�e�W
�d��9
�\6��0��0b�u�9�P�-!��z7�m�Рg
6���b���i	
?m�.Ǭ���ӈSۧ�[��u������>D=��!��+;�-��)S1����?�З#Y";Y#�C�c����z<(`a��w:JK�ɬ�l��jQ�$��[{Uo�z;�ɗ����v	�9�-Bg�+�t�����]��s+$��5	h�#���{�����U��Q���G��A��y���MO�Ox�R���M����en�	3L3�$��qK�\��JcC�j�"t.)�T�a��-A(�,ہ?�JbIl���4�P�)��q�Y?+ZpLX�*8ʃl�=�L�_�����Ehc=��Ψm��x@(J'p���DPo»�f웬y��\�`|�jK�!�;����(r��
���RO�&���&ݙfV�O�|�B��l&YH�h-(}��� ����m��	K�"�S'�o��pC�g��ƺT����4�m�%7�pZX�b�a�r�}%���6)��$i��%�!���D��w��ǁjҬ��.�C%~?8�lj�_�=�3i�F������*��{���8�%���}�aƃ�f� lR�[�����fAV�[����t��r�xY�0����d��O������'f�7:K6�]YL����k��0�O�k�2A�CiL�/������xgr����}�5�4|�{�>s���ЂC��Ȗ�	P�8oڅ1A�����OCl�.��<]}D��w<E؀�0��k=��^4d�T��DH׶�����S͸�	��P#K����C���a ����b�|���m�:D�IVH2���G���	}[ʺ9x_A^D��A�D`%��^�ŧۏ<��k�������1�
5�K�"���t�v��`I0����r�Op��uh���az�F �6K��N	b���g/,&��16��8����I^�b�iW0l��kC�<x�1��==��=4�l�MΊ�%��-�hG��	~�]�<�Jf����
������#I ���Y��d���&t��\hs"A����#wH��Oߒf��>��ۆY��v!2�ƴ�Շ�Ge�4yj��\V*�5����5��+$o�e�������!�`�E��=�HT�����S�6�r<����j0~k�͞U�81)Z�1��#�G�Ĥz��U���qt��~�	L��}$�A��Ugw�*�ܐ��H�+�1M��&h9V3Q�Dҷ��q��q잘[�R�>�{�}�5^k�����j��)�첉)�G$v ����ř�;�.9��Ȅ�106���㝩�Ц��jRf+��a���/o��>|�_����^���ׄ�e=�������WЁ�n�Auc��cë���M[=^7��ŉ��|����9���b~�$�.����jU���Pi�}Ĥd9#,ޯ&/ޔ!��HN��Y0��·@V��~���8��r?���߅ �Q�0̬��ߠ�>]���t�"��O
J���v&�,
�/��w.;��`S�7�3h��T�E{���J��/��Fp�?׬T7�sm�0[�QnQ`)�����\�~�v��f�T�7��ȟ�;�t�z!��X�c��4,^�S��-gf}�"JSC�t-d!��QQ1{�<�A���y�-�{	[�`�=B�P0��2\H���}6�v�j�Y&m��J��QL�V��n�6�C�|�,�p���V�-�Ty�������Y�j�PVR;��u3�<��O#{��MI�vR�P6B�j8
� X�J�O� �nу�t��r��+���_H�w)YQ�)i͢z�Q1<�d�G%�ט@GM�%�0߅YcJ��E��֣�ƶ�P���������琶p`:��bb(����]ϧ�xlՒ� ��p��U����;�ʥ��Em�C�:ԧ�� L�ks蜉 D�@��~��c�A���#��ˍޖ�+?���h�S��''U���+a8_�z��j��UD)K���&��k��_����Dڃ�6�����$�	�4�fP)��p��MaL-ӫ�N�f��W/xO��W�})���]�ۭ��C֕m̲fxh?�z q0����,�{���r����7B!�&9Kj�Uh-4��;��'M�P!]H��sjM?v�s�l�cu���0^XZ����a�++�GI.�͵���_�ğ�?��f�lY��
��e,��6��/�{�������S:�J���(����xt�V���h��T^�%/E��zG������;�)��f���Er@l
�}��&O���-��0�Kv��58���cA/g���w�X�	��j8]�]����?�Գ�5�Wl��y��/[���3��k]f�Xx��jD�]���{[<❽���W1`X�2do0��cgXghX�t�gj��9]�L1��R�D� )+����5ƑQ\�0wtz��L�#Jj���c���$�	��֐���!e����=:��p�d��Z����#}Q���:�s�y�]�������e}�Ȁx��)��&��9;�:��T��WE���ۚ�p������+ҟ!㕜@���Vy����6
�<-Nꆜe7�[�;Go��q�6�l��JekPG!m,�s�!�|��i(x�qX�'Q�㜟��ֈs3.�_Π��,�mc#��K�P	<��'��^�J�ٳ���iD��&t��v��"+N�M(q�w�Q�9#v��ol��.�1H���CiaH`�G�DK.�0���G���*�Y���!8����~�G��z^��c<���_ ]��գ-�2�yN9�&����
d��B�=T����l��bхM��P2��;"�Y�p{��c>5U8��t4��O1��-�C�>���f��0��e�m�9l�+��]/�ת;����<z�[�2K=���.�}G�4���t%�J�N*��
�̃�y���_+D~�sET��M��W�bY4��j�.(to�v�y����0�R�
bv:a?:}�f���K��2$���� �������3��@ݳT_'L|�C�+"'0A�~˛ce�P�~k�}�%�d��[c9��y�'�9�㪂o7��C�&�M/[�Kg�(�)��2���>S�&��a�/��]���jS��ۣ��3%̞W6'�A�7DQ�E-;�?*o��}P7����f�A�0]DT|U��\����& *�����8������O^��<Ւ1s�ׅ�ʀ�v�9�kQ`%�`H�_Q\@I��`$�GӰ:�D}C�-��m+�[T4��4��(0I<fM@��f~�o���3=�F�q3�K�(��"Xt}Pξ�ފ��Q;Y�1�����'|R7��A��:������	Q�L��FD��צ-q������ �,�����{%�1�ߑ���-;[�-�Z� _�i�9����-7��`���#a�4�-�;s7��w�h���I�����Vy8j�vHBG8E�u9��p����	��ӿ�c�1�N�4㠋�O��8��f�7,����$B��3��� ]�I|���3�|JY4D���NTk���&Ȭ�ߓ���:��	1@��?�ȧZF� ����*�b����W��۽('9��E���dEĐͺ�En�)~�:H����wn�M��*J�$V��?a���'@���O�!�9��Ef<�!�wr|ߙ����m�me7����\
A�����q<����K}����YV����"_��`#9��&p5������ϊ+a�}u���B��k(t��(X����¶68��R4�ɑ_xX5h���@��xP�^��U�\��G��(�F��Lg��&ԟW��������<*8�4?�k����[�l�3�l����9IE�=�L-�<�d5�r,�Dp�썘7�Զ�f�}�|m0�?^ kV�+�s1�3��B���U��|���iH�l����}T#{jk���gq3�ڄ�̜~$�D�yL��t���x�7��r0-����d�;���(��=�)��!ʎ��v�,�{*��F�a�`�t񂓟qde�Х�t�������z8w��y��,o�:�r^����O�@Twq&�`�w��-���;L^ϲ��J��=8���}�[�(էSG�����jJ�#ܘ; �`J���C�^�P�n2>gޫ.$쪶~V0��Dd<b�I<��]��`��0�+�~��.��B�/�䔹V^�բ5rf��=l��� *P�Z��Hv�,[#� �;d�҉�2�x�U�U�ʉ|U,J�mE�B��E ����'?�G���$_���5e���?{�ăK-������Dʲ�@�߹�3�Ꟃ<�	�ۨ��2�c�t�ge��k���lm�7!�&�Up�f(o�jc��IY��i5��Zhd�����
����;�g�X�4^�>���}{����v�Xj�s���1�s�6����e����N�K���Ѐ�fJ��r��>�G�#o�7�8OUD3q��vsxg��-�̩�r"kc튱Љ�d���{�����(�#@-T�}X�Z˗Tr�SV�vS��L@k��m`�����ĳ�(Gօ[rXP�wLַAc��ՃEԊ���r��8+?��y��So��y�H�XL�üܪRe�GG���F͠hT_%�?�Җ�7�e�޴�ke�
�/ĩ�֗�	����j�n�ѣ�,/:G��%��H�sN�hhG�@�{�˿i��7!K�f�2Bo�v��af��Z��5e��:)4�&I"`q�|�f/򐩝�Z�\�t�f��'`Ǩ�L�  5Z�ً:P�lέV���z�9V�P�u;�Q��*!=�"d.�@���"ׇ� �xQ5��hoꨟ�O�2Ь�z�n�cf�JwBn�_�==�M!"*�\c��7
�~@��^c�	��|�lsi��؆lc3C9����^�t�
ʿY|4��1�	䬿k��0�Y�� ����%Y{�w���ڥ+ �s��9���<>(ma!�/h���c��@_r��1�<J��y)n�4��Z;e�J�c�u���8vjMaM
����%���lF��)!���������^ �y]��+��q�8�c��V�93�r!0,��,�S�������e����GsKd�z�N2���	?�@'���}�
�L$��aҫ�5O=v��h�NV�g�N=���bnǻ��}q��F���pHo��7 �����3� ���x��z G^����a�+�5�I�m�%9����?��c�[8KFF�3%ãXG�n[�{�8h����
�&"h/����e�D��T����ܯ?�)X�	��H���t��&��aM�p'�Ӌ*P���0�ٶ�.Ո3�rH��Ԃ)��4x���C�`�y=G�f��sx�Xv�Th>%
2ϼ���G=���h3kv�}9�����o��Z�ٮ���݇�"#o���~i�~
l�ܤ������ӈJ�6�`����%���#�U.�f�-�f\�=�aF�Pj6�"���(W߰3@}LE�����HlYR������Lѐ�=�g�I�1%�<i)�X�i�>��$d�=t�R��P�WH+Lj�pҼޤ�"v�[pSe�>�\��tV��yX\w-�$ ����~렇V����A=�-�O���J&�21������D@5�{��r��kƂU
z8	9��,[�d.ԟ"��#�֣�-AϬq!��7��0����1�\�'޸��T40)p�ӻ3`:Ђ�R����U�w����Z���W漳���Xfy��v��}�HB_M�'����<ьπ�Z�a r/#�A�&�f^�R�Y�̛�{���0�0��Iuz�eeܷLN�伌\��^u��8ˏ�SW��,I�JZA�_�����<$���*rNj�W��v<�vΡT�S�vw	��V{JK ��'��2�^�[l�A!b���S����/ن����pBe��Yp
_���]u�V:������Q�1s  ��qd=�f�٥��m�&kE�w@ړu�0�8��!d޶�0�fWv!F�~pµ^u��8:��Ep����r=J��G�=�,F��²�C�FU~j�i�ib_�4lF�f8�9���Ep�
���Y�b��֊1{X�I��B���������J�ho��i���=[�ʁ-��x�Q�9����a�>:�iħJ��I�U|��"������G����W����w��AAd9%7a��1�8V��Ð0\��e�e�5�P��D0�!bl�4mT0%�wn�w.������V}�Ϫ���Vs���ӠrVw�$\�)wJd�<�� �"�o��C��!-P���1ϭ�Z�ER)w���������[yH("�5����kH�>� S�����{���Aq�wMl||3H����:�IR��A��S��XM���I��1Lm�r�T������w	t���-�����pm�s�k��+��4�C�62��FD�V���y>�0�A_oJ\�E�x[R��F�\��)sҫBw)���A����l��Π���2.0x��)����J�ω��J���P4����@�o�v��Jֿtk�TV��R]��ӵ���d(�*�^��É�:�5K����h%sF�҅NEٙ)�U3�>��X/�-��O݅���1�X�Bbe�mt�}��m*^��>ď��B�n��2[�*�L<ޑ��Â?ʟ^�=e6чs��Z|�h�6؊ͬ�r��h�h�,�jz�����zl"���?e�g��Rӷ4�Ⳛ,�����"o2�����[�+��9�x�keD�B��J�?&�W`t��#�0?<�`C�G�i�H�h&�f^9��N˃oG�a0h�"xr�*+��` sɓ8Fُj@����q�³�[����	|���XsƢ<7�� M��P�=��\c'�]�\���y
�v�6<�y�,]pj�Q@����^݅T�VF��m,!�Bz�W@.��`�rŷdDF	��.I�޿f1 ��9����L=e1�����Le�d��I��N�禴^�cͳ=6�Ϋ~�u��MN̟9��3�����:�VZ)���J�ӨH(���!T��ӹr�jE��<z�cS*�~�y(jc������s�������3-�R��p�@�o_\M��nuoY��w�J�i;`1�*��/�wP:�T	���1�\��{�0�dvE6M�4�xc��& S�	������u@���G(x��8���N�?Q0�0E"�e �v�T����ks�Oe\M��M)�3z�)���s�֮���X!������i��
��׏��Ѭm���'Ms�=���Q���i�O�U��A,�G�t(��m�b��I��o�tE,�|����fM1��9�o��K@ʀ��H`��߉LI�u*k�e�~._��A�'��� �A,41gw�=Rh0g<#�]��C�__��t��k.�Ha��0���,IDA�6#���m����M\/	��ǧD]>�^2�ޠ�f~#�\�j� ��Y� �&7 �KaU�d�՞2B�q�OD��ח �Q�00��R�ɩ��eS0��em�����Rҍ��V�X�p<�Q.�LP3q��2��J#�R �.��날�X܍�o�੥��'6Y��h ȷ�,��hR�|7Y0�PSx�����R�+��π7+lW��u�}�)�ɳ�U3SG݃\fh���r��P�����wD������7�-Yqg.n������;/2��sRɈ��n�=�4!�v�Q��=l@������Y%ƬX�휻�����s:���"�?�q��#��C%Z'�i���0���5F�l�_㕵��Ak�� ����
(ǽ��J͉@��5�i�6��t��Zr��eB�f��v"G�[
	`���n��Q
�tH���qv
��|�ep�g�4����� ���z$�~�^�W@E2 x��/�^���1SoD֙���-��H�'���]x�.���d���|X3��߷��#��o�t�ԡF�'9x�saX�+�)P�W��P���YXRr� �X�!L!P��3���Q>eF��ڬ�>Ojf#��M�7��s���U`��y+�>4���(:��Q,��F=6e�%�#���c٩�B�S ��e�� �9��mWmt�&�n�2� I�|,�V1!ǐ<e�lEnVB�i����zZ�9��`3u[��.�|t�cd��{�n\m
���ɯ)���^��Ef����Nbxd�ٛ���Z�6�6��`/��`E����I����|A���5�����V���4����ݙ��t��q/�(�
�ĀF��^�P�,+:[�k��p�*ա��">��Z�ю%�o�:^Ѓ�-J)7v�5D�`��o;�vp-0{��Q��!h������g�F��↉�e�iy �5��_Iʮ�@�������29��8y��e�<�\O�йSș�-Ԭt����5�e��zM��7ݘ((+A�t_���q	��~��.�&��K#��[����l����v�Qx�خ�js�q8��r�;`�Z���c\jׂ�M���#�e<[f�=�x��� �d@Lڷ4�1j�u��d
�_o�N_l7"��x�4~��K��;���xe������!LnoTw
��$(>�GG��e�]��g'�w@��2.
MY����)q��L�y���7�������rW�����o�ɘ�K���8��"�.=���*�+o��N1�#l�
:K���E.
Pe�U�1>���DF����:EF�O�u��|������OX.w�/����J�4�+TY�x�۔�S-&�c�6���L��j?�o�fA�>���,O���7XǙ��E�����1���m,S�sN^��8ωC�i�	���Y0�����ZX��y?%��th�Ff�_ZK�$�iA��]ƛ���.^dE7���m�2n���%�
�X�8�'��olF�CG�F��G4*�L�[�k���I�8�تމ*�+�@�[g,�c����^#5�
�\����Zg���hz~�����:@����~9e�v�T]!pV��E�43��\���T@�H}�BRe|;��Q�T�d����e]>���<�?&2?��Ť�h΀�Y�͸��K+�ݩ-��E㔇2�=�k�
U��0�yMA, ���s�8ذ�}����OMp���R�����jFg��^'a����ֺ$�Q"_;���ܘ�>`�:\�Qr{�=�^���Z�%��J^Zlv.�,�T�!X^C��F����UN7��6g�#L3�Jפ�H���[	.ֿ�^_ߜ�Z��C���_�hO�cX�u�m�H<B/ԝ�.5��2"~���!iu�&,��u��&��;b�tń���Fd*�}���]S��T��0m�I��}�:e��&'�q�ܠϚ+� �2K�J~����T|��|w�]�,�Co�y�M�Ί��|�}b��C���= >�-gq��2�j@���a �:W�p���.Zy�}t+K�u$$%�;2ڵ냉r�������׷��?�'f�G%R���\NR��tW]j�J4;���NZip�ykrzX_p�����[Qv2�,Y���1��@�.�F̚q��� _�pa��\���}��h�E��k���ם�|��g�3�z��^�/�T�:Y
���v^�"�)@����i���=��d�[HrD����E�
�n�r���2r/eO0�G 7^⦠*j���:Ǎ?K�����
�.6g�4sMi$��0��V*���2V	�;�"��/��R#Y�	.,|D��،p˰��%�}!�`�L�u�RE{��>�̥���}[�U�\Zc���v�g��ێ������Y�$�#*�5�-f�"�ȼ�:�l�%ڽЭ������`7��!�cW�H�9]\�'න������-�{�MX����ƥDC�/"��R����P�A�jz��Z��껟W����\<~�Ѥݯh99�Y	�
}.cp�$������;��R\�ƀM�`�V�gq@X)�5_��/��ә�*����7Ci~��,��qFN�_������x�{P=��t�d��3��
H�|��Qt�y1��(���]��.v��j�0�-J#WV ���$]s�G[��9M�j;��ʆGR�;qC�.B�Eb���Dʲ��bv/�����܍�����M��`�ɸ��?���$�0��(AA�5\Al�0��#g�Oy���q'>��'�m�'�N�{�XI��Ք�%����~3L4�l�w�(����@�cp��`���Z��ůѰQ�#��a�����H�'w��؃����w��(@*�{��(���Q7W5�0|I)�I��@���zB�>e�YҾC�����腋�Ro��]��Jg��B�<KR�<`v*M��,>kh��&��'�m�E�~nF, v!�ˬo���w��T=sH�	���'�2,���;�PVA�KGDi��r*(�%zu����޳��.����M�T��s�� ,���e�_;�=�3]�=�w��_9Pqui��X���1^Z����+h}�(+���$��T�i�ݶ|K�б6P��=�w h��0��XO��?���\�T�0���}�m�g��s�V�=��3\i���g\V��L%���|���"����������`2���Ū��v��ؔ��
O����A������QN�$t*&�PQ�1N�_0'0���ӱ��vA�u�0��%�g;���L�?a�I�hl�6��j" '��]�ׯ9�;q&����.}M��=O��g�� ���^�ǓF	�(��}�#U�ժOe�WyZ7��몕&�LU |n�>q��ўi��p�)��H��c��u���o�O��o����S���ś�6j����PN�.���Ys�kU����3n-�����ޜ*½�^3t.Y����>�2�V�p���W$�#`���H��xP����BL�x�l��iq�y9�ԝ�~����cԋ������?��z!S̔\h�r���4��*���1Zһ��ʥ�L��Izr>d�q�tXhB-�/��V�5�!ak0�E�^\�h��Fiļ����>r�tV�������d��Z[��ݱ�ِ	pL�m�a(k�6�����0�#Z�Z��Bf�GǗ~���W���gaO�S]!Q�_&қ, ꨼w���ܭ��m:x��vRq~��XA��4�T������q�ϕ�V�j�l"�wh����}���,}{Gjo��y����rg�� �G�S����T�^$OoN� fv`�,��c��A\���<�@Ǵ_�>Qa��&�s�5I
H�h��r�lSo]#+#�lqQ��D-�c���C�I=�+M�>j>�=_�Np��qܚVa�nlE/���VӚ������z1�5��i �Z_�漼����zJ2�0��[�<�J�|�*���H����ź��5��	|�3ٵ*@�3	5�vF :���Hj)-SpvP}`�~�h��?���!�ݱ�E�.�](��)el�x�=��v0���m�0H.	��{Je�������V�c�3a�i������\�Ta�-�Ȅ�-�"�>���҆A�dZY�S��<���;FL���<8�D�_ٵsb�_a�!�2�m[i*�(o���t��^��?���0],|;�0�N�}���2Mګ� �^�Y_w3K���bj	;�燂�Q��%�l��	��pX�Z �����	G}��x��fZ_{g��k���{�K�*�z�9!8v���]�+�b
�Iah ��
��z#�B1�&<��;��!��duN)��#Ϛj� ��̣�^φ֦Q�wCIR��n�8���̓a;M��G�znP�� ��ۙ���-��A�4�%V�[O%�v�K�[@`"7H1��!��Q|��I=�z,��(\y��l����gg\O]�yְ��+�����Gt*��#-��t̓������M��>��m��L��YȖ����M����w��t��:5�q�Lw��� �ێ�A=T����hR}X�]Q�i,}t$ғ�l��i*�rC.���٪��6O��b�H�������!ǲ�Ip�5w#t�W��9u�?�����]x����"F-�����\g��g��BcZI'���Z�޹zVz"�m�JƟ៣@�����IY����!�ܖ�@��@�,9���	)�^�U�$^F�X�1��,M
�L�����p@��2��q�h�	ӂ��i���x�]U�X)��<���n�]1�!��*��wK���m���^WGό�;����������E�l���mw�SsC�Y���A�7@Z�23��2ʈ>F����5��|y��$�_� tQ����x���R�ڴ�У��\��#v#�X��z�{_��(��g��	�;c�Ro�	E��l�O���mi<�Q���$�V�r�x�'�I�0��)�A����3J�{�t����7����v�c�V����p3��8}����@����	8pc�D�K�	s]9IA?~a�I�lE*�h;��xg>7g�:���H����_��i�z<(����?YE������tT_������M͓��4�N'`�OA�C�˔�YbUY-� ��Ѱ�"���ՉE!;�"Z�З�����t%i�nSZ����4�ݟ��G��l��&����.*L;�Z��f^4r�|ʓ��&�CsX[C�z�����Ι���c%k 򦲽�)�|�?3�q٢��&�?����y��Q�0 a)��܏��fvl�����<A�P�{���y��:�S����;�LL/�ؗ��;v��.��Z�&䀘�t����"��`^�����YQ�*�X�(�s3\�yГ��1���r��2��-hcI��5|)\���g-x~7X�Q�	:p�,/�LTi7)����b��h�X zpNڏ�e�&��zM
$�f�O�J%VC�v����I���	�`0���G�M���ԯH�v�"�Q�eޛ�"�̕���|�d�b-����7�N����p�=#��;�AҚ�3~hR�Vz=,÷���(�=ci���l���U�y��(��՜�o%�3lnb�P�����zJ�>��]�Ͳ����W���$D�S0n�Bm��W�\l���������WZM��P��#�������y�++��ک�N�������pa�yI�-lg?�E��SΜn$�cHZ�%YV�l��+0|��T>��;��!/�?��4�ۉ��#��&V "���Eۣt���]й1~6>O��c��H}7�u���z4��0�N��$#=̿ś�R
�J5�wY��-��)�cױR��q����CJT�B���@t�$܌e�|�"�6�N��ȋY��&������)�+�騒�\ճ[J�j�����G��q�A�'^���<��ϰ*Qؕ,���*�b?&�h��t8�Sӯ�O�2�ً�6�(ճ�P�-T7��0|�>��<�O=\��=��Rq��Z�c�����-Ҁ�����Ft:ș�I��N�)�D%�3�93�%W6@�Y��&	Wm˸���A���z�Y1I����&!9����>�	���?=`�髷)1dx����1���)���f���E�����2h��E�����OKe?~���X�,644p�����ڳ簁>:?r2���f��q_Ǜ l������BSR��"J��{f�V���gv�K4���ObqO9�����Jt2��g\��G�%ƣ�\�`�쓧�m�+�NsI
�-8 e v�BB"]1_o=�̘4<��|�3!ߢKa�����I�Ҝ��z�2B�=�5�s"f�mO����eaq&(�Ս�@#�������_���C��hL��<a膝1w���5:§����\u�����@[1t֔�l��jI�аX;W=@���-P���:���7�����mw���貇@p>��>�+"�v�������<Kcho���z��"�c u�JU���$���O�X�NQߒ���v��-��E��'ldB����۴�|<!q��>���@���CS����>��3^(Q�?ÌQiRD�Hq^���P2�6�n��-0�z�����1wWAUFKC�[���=�*��O0�n;�r1��\1C9Y_�����/u�����3�2�����s�HU�db�G��Tq�*8��w_j>��iM��k����wa�>����j�(�����lo��\�e�C��گ���*�56cu$��+ /�>CI���P��]M.�
���-h�������Q/ �͆vroE�����e�
o��4��E��=�XB-������W�v����A�|�R�qn4�ta���w2����7� ����չ6�Ex�+HX���^�TL�h�D$�m$�st��mPV?Im��П�d�lU.� +ԍ�oW�	Z�	��&P@�c��������pm¥6q�a��@o(�	�v<��b�G������[1�y{*GTOo��jd"/����"�0D٠ ��+����K�Бb�Ō�@��O�j[|l��/��7or���R�N ��-#�8��<��^�,T�y� (�T���y(z��	�(lVI~�"!9��YU�D�f��ж30�U�eF�SGH�e+�`�ߔ�@Xz90�݀y-�yINpJݷ>J�սFh�{Q��1�_��`���	����%�k�[�g�>�E��M���
>h�^�T�*B�	��x��(�O፞x�,��u.��j�H��.BI�g���V�j����4Z��q�-�sN*�1ɥ� ϩ�L��Y�ζ��V��BR�XT�����X�t�������h.h�M��uQ/[9A���\�ݍF��\矑�PM�Lw�ֹ=a�$��׀�"�o�������K?�@�c;V��z^G�Ϸ)�����pנ� �Low���D�G�sy����4��#�
�s�x)���O�I�=�QN����&�9���Y�1�y��e� VE�&Hq&	�&���2C�j�5^���T���*`�.�5{�K��v��g\���[��giƽ�0!.��ӳ.ʋm|�OŢӑ��Zj冖�.���0W����)*_�N�? ����`s���|8n��͕��t���M���$^�3o�Fz�|y�SY�f;�Z�^Q�K�FP �k�dg�6��i�1W�ń�t�[�=��if�S��*SW�܀���V���wTF>u�߮�F*ĺ_����6��AO�2�������(XUu���5�B���Nr��6#���!4������SqDAZ�0�Ip�9��!�M��N~���w�bL��ًThE��1aE#C1'��nz���-��K�!'|�J��%Ir����
�- ̤|��	�h�z�zY~���B�>���$G�l��ąR_��
$��X'M( �_�[�B=&��Z
�B}�1~D�
J7�DL`��i���hXB|�+��Nx2ǋ��%�~�ym��v�l^��B���jv@�e�]��~!���g^J_X�^�1EiE���Q�����u�y�Ξ����ۥ#b�����8]?��d5�AI�t@�e2c&P��x��G��T,��ܨ�N�Eu8�������2 �����̴�&�I�4��5Om\ x�3ò��]l@��~/6�o	��F�hev��0��鏥�]1;Xi%Sw+l�{Z�JH����,-�Rg�݅My�x����椬��*K>�%��F�����
W�}J�o��	�ħ ;x˰=�_�\x�`�@�H��Y�b#{�݇�zIn+6��k�L�H���<g���ů�l�E劌)��;m���@H\�v����S�q�9��rE�M�X�xPn�S��O~V����ͤP?w�p����w�:�њ8Tj{eMW/�0���dq�K�薮����������s	.�r�vú��@u�KY�?,��o\�nھ�:߰^�u}E�S�ᙦfKa�Nש૑���,LE)c��L����z�4��Q&�r~��@��^�p.�x����W�8�ַD�)�xlF:6�@ܸ{5$}��E�6ȭ=ecy�����m@��&���߂\!E9��>�4��V 
�9�t#:��Nu�YLY���bM�vP1&p��%T@�����d�d�/u��7�A���K$�8vl�$�L+Ni�*��&���ҕC��o�ޓU�"�B��猫�|�}��'G����Cs�$ �琗��Nt���Fi �;�&9aՐ��Nͨ�J���z���B���v �2��_L]xg�E?E(�˃���B�x�J�+�Ky��H'��@E����-	���M��k���c�t�w�P����t��]�N�k;����!|=�FI_=�>W�Cr�"�}����l��-��N���O[�#WPMS%A�o�}[��U�+�]U�Py����u��Ղ:�Ŝz�J�JQ�G���5��zdt��Ar�z�_B�!ˈ�1���(�i}g�a�t�&
^|~�'��-���V?���ѓ�����\�l�Ѫ�}�i|�cI�i�	�Vܟ.�0g��~�ׇU?-�D8EP_2a�:"`$h�ZbKNe���m#�y6 ���$$7Q����H�^��QL�,�y"ĊZ��e�'°+��B�Q�|�X}̸}�cG&�ű2xf��da�f�jF�Y}	�˖���JT�ԋ,[R�uJ�$#F��r���6wʩ2�#g��1�Jc�K�*���5MOm�����E�����R�/��D�{�hEKS ���0�ޱ1#��߀��ײ0�_����T�#l�Q\���bY��'%X�K*�׉��p˱�S<�T��9�P�_V��^��
-�,V�7�P�A�Q,����6���"�k4	�3H�
Ih����GM�G���G� �����3�TѼ��[͚�=��!�x�%�'Mo���M)���Y��9�ᅜ�q 寘���/��y-K�~7����6�6�]9��E���%}KA�Z��T�S
7��g��p�b�R�]�R��Z+|�'��eY���z�c�<�9�N�if"�x]��2�ˀ|֘V!�@uT�aJ��Y`N�}���`G�{������#x�KjE�J���ђH�tn6�/�ö�Kv�2b��I�B�/��_�;fnq��^n&˨�n��������2��[#����%u����u�obd-W>w&�N,\�x�l�:������ڗ���𓔷������pj�����YI�����E���g�^���f���"�P_�	)L��ר��������;��pf�J�~#��O/�Fn��R�-�l7��zL�tCC�H�uʨj�,������������U�P�5��M�7��ݳ��'�^�����嘷�����7%�/��C<ϧn�9e�1*;�>K�$+�t0k���_y.|/�"k�6#�W6i���ŕ4����۵��s��]�"}w7c�n��0"��=�c.TU���o�	.�g�}pr���h���37��s�ߑi�iԪ-,�l;���U��<W/D|%��?��"�I�5�Q� ��4�h�Y#�H"�_8W��Ju?ˉ]vp��M#�&y���m�II-�w��;x���QZ�@M{��u5�5�=p����3U��a�^�O�,ŶC�I\����_�I!U|�4䑇�q)4����{_���2'	�"?7�
�m��R�0�Y��,+��Q��zQC4t�%�I�W,|-�v��	�р���N��m��L� ���i�F
�[$���s`�z�\�9�p3�2e��ձ{�+CtQ䐵[��=u=i^g�;�,g�"�"���>J}��-S��;L�$�\���Ϙ9%�J-B;ӑ��m���ی��J%����<��k���GP@�u��q��כ��&��	�ϓ�@}����+oe��ߕZ%1�+�ѽ��H��Ax�`//>���E���%�H�ȗ~@�L��������+�yK�oĸ��3�2�����w�k�2��,WCj��(�B4�ٚ��m����r7��`����،S������^iۦ*�0�n���V�+�"5�37s�CG('d���Ʉ�_��|��gI�:�y)����G0	����neiYwN2e�9�](�ʨ-��(],�N��xM�~�k<@quo��#2��C��P��̒���y.(8��Qc��� Q3����pI"�Ź�"����~�$ЈiQ]�4��Ӷc�v!�Nz��U�V(�l��|f�(� ���t*/TYLo�=i��H.�9D������iM�1�W�s�Q�?"'� }�k�Q��Guzi|�g3բ��!}�ܿ�t�/�U)�>�e�ی9�n��)��DÑ��A��Mn�cC2�`N�B4+��� $�1��雯^�DʋQ)J�{�� ���v�y�� b@}�\a�A@�;i��]�F>��DV:�"���zI)vǙrC��Yf9i ������j��_7�AAQ9Cn-�*m4(�_�Dh�,���wh�h��QP
q*���Z�\>��%���cR����I3�RqO�����[ڟ�;!���}?������j�s��^ûG���7Ţ�r���vv�N����L��53Xm�&�����W�`�w�n�����d�U����q*?@]��3IW'|�3�%)���v�	�=�ڔ�[^�ۅ������ �U���C�$��y0dԒW�31'p.���TaכCr�aq<�L������tg�ɰ���.i7Ϳ-�:��(�?��n)�_
� Q���$���q� �V^G��Cj�E�:-c�u�ؾ]�_9��H�2�}G�i�*D�ԦC���s��Qt�XB?��ۗy�P�)-��;�ŧT[̬??t"�
 �U������
�� �,��$�PA��`�Z�����Q.oϘ�I�)'c�GK���w*���5IaRc�O�ږ�24���0|��1l!b����<�?]���6��Ύ�k�پV���b���0|��٠.Dwv�j����o+���!�!c�ൺ�tVq�U��Q��}R�P�޻��u��_�z�9�&2 #m��V�~��0�Ǵ�4;�ؒ䊭��|�m�҈�<٠��#�8�����w{�2��3��>����B.�KM��>b�/��0^��Mc�Ϸ�א神%��vԑ��c@���~���H]��q�O���Sj������d�g����oWÌ$��̹nt�0�"�Ɗ\�w�b�
3x�Fn4��2V��O`M�Ӎ�.�~�_�����(\l0ss�iL��p6��Ti���b�i�lNg��bY��?M���ct��nO�ZX���5H�}�-Ȱ���n9*ݛ8K����<�>��� �p��_$��m�5	���xuy;��t���SǱ�9��x�-L����<~������C}I��Ӛ�n{�Ҝz�l-Ѿ�{��o��B7��ng�~��BÄ��#�SXs�9��)_[��S����ۦ^�ޱ	]������i���,�p��4uVǪ��-��oM礘��QV�n�Z ��/-_F:p�bz�u�3�rۑ�@��{��V0=U��֢ÓH�f�>5,=���w�mr�)���*C�/�]pxgy[�0�ʤ xT�+ �G�񯪺D+�D)'�B�En5M��ઉ�?��C����������\��/�s\_"t��&�`��|�K����?�����~1�Eo��|���5�2�0�x�e����19%���yrؘih�^R!�(��,�������|rP��q��|ܦ���B�����9��T�
n0� Zz)���C�eG���Xn(i+��xզ�uSWsҿ-���´5K� xm)���G8&�":iQ��~�����,h�̦0�v[:d��v���Uh�dNIBr:'s/�F�mg��ׂC���_�f��4B�W�M|V�k
x��d8qa����!�{���M�����F�!�����訒���D����ZZ���J$�$˓x{i��Ҵ ,�~ �����{���I���Ћkc�"+|V��H���:���/�6�Ɋh)�@���B��k���J��@\��;Uo�lD� d��k�fb��-�p=�߱���WWb�[�7�dNNr!��] �'I�c�������͂��|[3�~s�\[�B�w��+�T���tv�����(�I/��Zm��"Ȳ���4�ϖ�p��3Q^��Mת���')���7z-�M���V����DǺH�,{�;�o��wWn�����(����8ן�i?z���7�'�$���wF��a��]E7ɧ�'&t��:%�Ǩ����V5���e���t�U���l��:�h�Ǫs�ۿO����:�ÇE>ׁ	�^N�_s�x@��5�������+��o�˿���԰4�6�+8G1;��6���F��j>�4F#����n?{wc�?��rΝ�r��q��a�)a��+yll�g^��/��I8|����<b���Zl���q�P)a�W���M�c��ž�R���w,~*�#F�v�B^�r׃t�Nb�x���0 ���ĦHnqY��i���4F����>�Px��{U�@ِ�0�18����d\��7��ɍ^��V��H�3�m��f�d燈� ��7�%��J����8���0��uӧ�-����	ڗ��	?�%����6����~2��R�n�y�� +"����o܄�F��c@��	��%�ۓз�6(�z��I�OC&!j��(�Q}���%��fQ�v\�_��a4΅���������%P��6{�MjO�A,i�J��ļU������7����4߳i{N�~�l�b#�i{���g���j`j���'�(�!C]�(ݤɝYO+j�P�K; ���l�YR��~;=�d�V-�X�N���̛/13l,5g��������b<��G���:�@�4��SH�"a�F��E����� 
�uv�}�o�_bÇ�����nc�9�A��.%�D5�|'Ժ4�	�q]}!����S��!�ވ�����t�;�U�$Kİ�^�A�Ǒ��@��x$	���I�;魒,�z��}�r�n����80˘�B�����x��,�� �+B��%���=��v�"Q���J==h�e�C�bQ��^]�y�v���^R٩���eN�l��[���eD�P�`�C��bk�5�%�9����P����|
��r�&��|0��Eb�[f�.�]�Ka�:!F;~�B��x\��ڷ�W�YW�2^�>� .Z��S��}�{�u�Gr�� B6u�1��o���*��U�ߚhU���]�����i3���Y�F{��L�B�Ǌ��#��:���)®p��Z3ط)�~���z����v���+�iS7h)(�,�a��&��%}շ����,��:�RrZ�C�saf���-+v0Z14�46�}���A�0��w�~���lnሷ,Z������P	i�I�m�w}�U<pB�U�x6�*t�MN�if�C��W������B�J�%�*؈Ґ���!�p	r�40�*�N��Do�E?rG�[�@�7p�ݮ���XdK�o���D�Vj�_���[�U#4����2�}�YJ rX`d���N������B�ے5
y�D�9��r�w��稿�����t�z��@��q���7���jE&|a�=����X�����9\�G8r<GO�L;�K�RD5h�k:s ��d@t��N\���S��e^����ܒ��E�p�_pO)�F��x�t���m�푿��'���僇�<s��,�003�D���7
�n;ׄBH8���!Įf4L/���(# ���d�x�#��O����_�6z;��R#�N�mŤZb��uh���:��09�I4DJ
'_�9HkZ�,#^>-�g�t�CЀ���}�~Y�]��c����Ӯ��o{��'F����}����\��?N�=�vyy�d�{�����\� �oo G�Sj�?�3A��7�G1$5�ec���TCk�� A����4��K.�!�6J���\�� �������Q�h���D#M��j�}��[v���N5��T��3����dXo�������W-Wm�65DꁏT���d��$��������q�9�.�3J��lI��"�oKd#~�0�#ӹ�>xM���Kt����/sb�1K��B4O�aS�s}�堒���^i�V�fDP$��'����s��L��ׅ�	�%����vt�j��5��W����Cu�dpE��	�L	"-����-.���R�[#����PR������j\�����WV�@�<�Ҟ=�=��[����~gp%_ ��/�B[���G���K��z�����+��p���JKW��鐻�+�0���@���K�� [��9)����k@u4��	�����k��`Â�����,����	`�7RZ9�!�sKZ!(L����l�}$��T�c}H���<��n���a[F��DpCU��W�;2��[gĸ�+l�/���R��P}N�a���3Ǭ˞� �j�Lhu��5Z=fZ{/�����'K,Ǔ�
Rξġ�ĳ
y����4�~v���E��ƥb+�R��,���c�}6v&����=�̕�4�>��]���C�F��gG&��2]��R�+J$�f�R�	�m��.�z��=/G��1���#gU�$xe��хz �~fSR�ܶ��9�,��x'�KU�zL]���p�E��u#��eZ"�u��}s��w WZ����c�֞�5�J�@�%���\;�t�/�<D���;��%��H���5��;�*=�D�YO�#nO�ke4���AL�4���N�j�,H���8_n�4���H!Y�6�Ӱd�@+6�s���f]�y�\�����S?�#��X �w���P��*L�*�p�-p@�;q���ևՊ�'����}&;v�����2Fv��µ���i�I�p�����sD���������{{���*bJF#�u
��M���+��\l"`غ`ho�k�Of�۝�l��T;�Cz��u����[d�Mm��x0�_alߨ�mWvܴGz��d��VνEDF��|�� ͵��3��8��
������s-��>�@Q4Ŭ?�FYP,��J�P�,X�Ƙ=_dq4�55��+).L#Y]yn��L�"=��[gM�z�8��0Ǟu�(?с&��3��ٽ3���prR	�j�펹����>/�z�6�c���bo����9����c�ث�{�v�o�	�p�-@g�3��1"��)Bt��bb#5��vk�<����<&�~�mK�C��P�؀aRd1�Օz)�A�sŕ�,S�h/�W����5�3��V�qZ-�u٠�����m���b�_?�d�h	���w$9�V�s[�]O��VVK4�8@�� �j�X�h����2�ln]J<�#��
:�X�����W�k�.�������`q[4������yOv��m�l������UK��c%6����a��XR�r�`F>�U�n��kL?J�RJǝ�Y�#O���X"������4��e6�5��I�@�ԣ�=�h��ɚJ���+�4�����8��%�&����!�ȝ:_,鎸���~7=(��7%M^�h�{�����\c�o�U�ɳ�˗���q��t����D_�a	~C���m�5`��Q���\D�lJr�T�o!{N:��e>��D��b0�`�����󱂫Y��Cބ�%��JsU����AAX�{+҇u�ʋ��,�U�x�)���{�1�U�Bq�<(��� ����;�t�Wf���C��S]�1q�
��e�a�\��b	��üa1���%���6�b�5��`R���_�E�x�,��V�9<����Y����2_���>!| ��a�,��D�����9�v�H�ޔ����b�g��bhS;�H���Z����ւu_z���6`)����=�E��Ͳ�ߕeR�E��31�8���NbC������P�o��%���͸��>Qf�IB�{�pF�����l��@�d�����n:vJF��z�5¤��A���]��e"�s��zE�&�(*�UЛ�����]r��QN�sK�SX9�ܮW8��H����]u��6Е��V��.K���1�9��y��[h9�JClԢ�w L�nܖT"���Vz�1�4�#�Zo�#�/�ݯ
뚘my���j��Ϻ��F�^��F���!�Թ^JX>1Sʶ�A���^���}�
9���M��Xʖ��OpP���^ ��&'r�X��<�sr!�� ��a/��:}>�^&#�#S��z �rH�GI
r���=��h_���ž[k��nR�+��"�1h>�3�]��\��β����ֲ�� �'�	��4��Y������<l��P�j����
�3��g8�Q�S]�;U?��o?C�UՍ���?0���⥃7�����RT�6bw�r�G�x�r����] �y���J�c����b�]K��W��b���u]�q�k��ed��N1.)��eO��x��:, &NDVzu�O���cIp��ͣ��`;�,mhi�*I��gQj)���]~/���&��e|%5�P(�W ���k*�>�5�Q_Al;%�NB�����I��l)jl��(���m���*��qL(+V�7S��^o�g9Q��"�s|TX���&�����b����=�߻��t9���%^k��!3%*<��P��.��m�x���З75��9��e{e;���,�<44
�}+X�{���\�W���
.^ě��sc�uX&|���������sx����c^ܖR��E&舞͆x�n�/}֭��wi���ǅF�H�*��M��k;��
9wlCp4�X����<《Z�$�I ��W�_��ȍ,%Uǽ��07�R '���ݛ� 1Cr��V)w:�_�����u�������%�i�QV�6[�����b��C�M�N4�dٙhK���*�;�@9wt � Hm�R'M�?���E�Y��)�z<v@��6* �ݧ쩘{��N�T��g�j�5�Ӹ���x2�����6�J�u��d<UJY?���p�S�$`i�����`������T��5)�w-˼�}LFAPY�Z=Ϟd��V*�QAUj��l��8�{�ᣔV�t���U�b�Y:��PHMJ$��N�~_�$�hWF/��l���ڔ�YH��G}�J6/x���$nt�@�8������� *b40�lp�n�f�JЇH�	Ƚn�	[,�w�D�fʩ���z����R�j����j��* �o:�C9����¾ƺ!����C0�lm�#�������$;IJ�
kS����)�ZCC��2��_��t,�Yҵ������@��_'�(j�@�
�/FK��ܢY�0ѳ.���R
��t�۹�;�lX�4�"fjN�����+���`?����f��C�Fn�rV	4"��6w���鐲���3�u4頩_��Q�!�s��kp8M^ame<�)�U��	����xIr-�n���IAq_h�L,,��?��ʲX��d�����Mߥ9�m�X�:��*�@������+�U���H}�=��l���q�M��ïP)`�^�Y7�ֿ@�[}��3!8��gD�Bo�z����@����§L��|���m���[�)�;S%g%�;�2���s
܇�s��������w�y�V�����#�d��{�������{T� �XZ��S;ZMk�^E��:���������_�Y�Xnu;Yb���~�m)�g�Յ4p�h��Σ���O��8�tXEW������+�. �/�	D]*6�����a�W�:��c��2���+-q$���O�B���!rs�xx W��$9�i����K�}b���O9p]52�nn�5m�������[����q��8�Fk���֥��>>�(����P�2ů��ƙ?��X���4*���@"n'Vj����˞��~��!���m�"��^m�� �x��gJi�[rdy�n-�ؕP�x��uu�� ��慃����(���h�(L�VVc����$�B�o�s7%E}SI�,@B�{Z%`Y��g��*b���n��^zU=� ひG;����%��4u���k�<S]�&ˠ�J��c���1\�`�#�eL�ľ���f)ti��t��E�e�E�NI�Tw2�
�@8ڙ�M߯���?�k9��t~��o��{!
���������fS��HD��J����7l[F.�F�+2R7o��pp��f_�qw��Y��+���".bG"#c�֖3�j'`��@DƉ�m��T�҃Q����
R��E�`��؄����Ǘ��<�~r���V'���	k� �+K2T�W�O�If|A�Rs-Zr�'*��t�ۉ"���P�6�!^���\��r�;#�jZ�eۖ�.#<֬��f��r�:,}C���B������ֲ�+��=W�L�c������b�ʙ`�Cc&�G���{/�^�tN;���d��:k�]k���|3ֻ�U� o\N ���1��Y%��Q8�Y�%��J܍b�Ɣ�s;N�<���=��|�U+��^{ҥ�|q�s�M��*������_8ȱYvH�4LJ��`d���1O�i�0�+H������ 8����]3�x�*~W��Cj�-Ƨ��P�g�|�M�gyӨ�W�M��/G[�YV�G�Iq0���7�7��@I�:�뫚��Σ���o��� a�4�W� IΆ,�66� CF#�39
�p�*����Ldԃr�7V�"U�<��{/ILw��j�(�eA��/���Q&�n6�z�pA�q�2����""1�56iZXI��w"���&SҸ���eQ�X�H}�~\Z-�Li Ɨ�S������މ��7phY���IOѼq��{�]:�zͥ3�S����R�G���=?r}��O�6�Z&�m�� ��7m�w��f���*��H�n�Ṳdu�X"MŁ?���U"~N{�� C^�
r�i</�w��������3mr��f���G�\�vЂ\dr�6���e�B�GPB�[?b�t��5�pu�mI��CX��7m,�z�Vg{� p���
�5�W|P��ng'ѥ�֤��~�-?�@a�x*��s��w�%��B�m�0�r�v�b��J�>s�jEN�ޘ���1�2��v�[��;�Pn���.��rX;;ݪ['�/$p����^B=Ə\|�P�Q�`��Ia�K�����9�z��w\ Qj��_���zTܻR��!�n"�BT��T��O�xf���eYNC�{yuX�'M�#��E+:;��ޔ���f���W;ZЉ��R����S�kBt�i����[1Q.> E�5�3�7���t�鰝���b�Z����&'W/��n�s������_+ٮ"M�Ӫ��4�uH���iT�4�܎���@ȥ� �~Y�`C���y`*Vn��������*��l�$�ښwj�D <���KDf�z;T��T+�U�v^	,>�����"����#^�I�mF$��/w$�V�lMd�aI���N-߀�(Lkw�ݓ�4~JY3`�hSo2�}
���%�j��b���܀(?j�[6X�s%��۞��)���ȣ޸����;,���s#�c����||�<��(��<�~i���h࠰�~m�"��]h�_=j}l8����.�[��I�ZЋ~���}�ط���!B�y&�n�dj��$ߗ�åMrT|0;����Z�Q/r籭4+\i���V��ᨩ�m���[c�K5��g���:5֖�d�o��7����n��O>��j�^�c�w�(�P[���V��J�?��
@��9��ڏ5p��D�8�Ty�}]v�����K�ebׅ8�Y*�Br	^΢S,|Nn�ܹ]>�����w�����ZS���>�S���FA;�$��nHP����(���Z�!Q��	5!"&�)��
4���(��/w���2;����"��S垬M�����ƴ�ļhط2ݗ��埆�a;'P+a�5��:�m�IL�u&��SG�8"ņ�m����y�ߗ�C1*KHϻg"�{�;d��]�\VQ+��2�!ی�ϝ$��)ٮ7[w�CN<�V����=O���[��$�V0N��M�����sJH�iN�9R��K��O�\��L_-���O�N|��k�`� 3:�� gێ����ϲ��Ү�*+R��֜��Pʀ��J%����(�l��^�;�w���p�
�仫"_m;M���������kw���a��~������ռ�Rه��2��I��Kv�q���P\��":Z'p�#S<��l6w'-���������2����ߺh*�9(Y�Nc���f[!�{�t�c�*`4�)T��di�(V0�9#ʸy�k�:�B#�	6n�����\j%_�8P&��[���.��\Y��m�Hc�w����-�r��xΒ�w#�qUƅ�r��@��)�P�%-]� �6�;��~�ֿ̒�������Y�\q*��&�ت��|Zg-q`��
[+ �a3+�d� g����iv�����`�4"�fQ�E��i3�2���C0M�bp���&���H1Q8L-�+ \��(5����8��ef��WX|5�}- ����Ť^Dxx�B�*{Q�v��%"��V\���m<�pE����r�1�W����vq"j����5|XVWJG��5�G�Џ4��[wE8{�,P��b��u9����(<�̉50��1*���=@��lfa��z�!*��Zk!����*A����%a��`El�a1�*f-1��f��c?@k��M{��1U�)[�Rk��>�]dІ^w�($p�8��U�K@B�q��,(z����!�!%�1ڔ����򸍍(�e�zfx����k���	
����Sx�@
p��C��5��V���v��p1SBѨ�J����⽧�H"'�iլ}�nȓ�o�l,`h�k@;�	I����[S�EދJ�)�h�ΟQ�.<�����?��u�@f��,���E�.���  �O� �HPiϞ�;)�3�1y�.�{'Y؀k
�'­�ګ���t�J��}��\܅4Kz����(a"��>���Go����w��`�t�s1}v�c���F<�A��%s�C/	��7/o��2����6���%���������e�O�Wb�s׳?ťF�c*S���=��l�y<Tg�9�F['�4�jZJ*v��N�N�3��2ǬG�֧6hb/�9,�f��8����v�tU.z�,��/�Ho��	�r��\h���� ��xgN���B,	C&I2߼����'D�ݩ�O�2ɛ<1��h����� ��
]�G��:~��U����"ڟ3�X��Tށ�B}���� ȑJ���-G���s�V,�w+����Qh)�7���c,T����1�6B�z�s��oe�A�N���u�v�`G���&A}�8K���1��O0Z�S�Ԡ��G�Ϣ]d�>�C��j��EՃ���� �{I��e4�5Brxӝ|�E�Ȑ����Z���p�����;@w[��{�Z��&]��S����;R�Յ�ro��V_ʕ�� �0��X��Ah2��:���.�`Q�&�d����X2Fl��7�K��EK���֕6��U�!n]���X��՞ڐbsv��H-��H��i<~U����'��^_e���@�J�@�ܢ�f�ā�j_\��1#�J�����D��"�o��߱��Z���P�w��28�����'���=�F�QJ�s��k,~̰Ѹ@=� ~Q$(�&A
�����ߤ�}[�����Bq��h�G��K^g�8�t�r���*���1� \�T�S�H�-���T>�f���.R3��Ýڃ��<p����� �
;���å=Rυ��9�p̞�'��p�X/CG*=!��e@YB0� O]��!k�#�/�@_���`f��	F��|yyW������M��I<�G>�6�4���9�'�W�?ެ�7��{*�8�Lä��4����i�z&ܗG������dt��8���oI�x�5�/�|��"����_��Ü|
�$���Z�O-(�n孤k䓃�b�*�k�X�����i���b�$�qV18Ȋ�
Z�(��=��7'��k8�H)����\p�d�������I���k����3���87���B�#Nv�wh�)f(d�I��p<Y�kK�k�=)���4Q<����:��C`44+�PU/��`$�G�G�����D%5��Bƪ?!_�}v׮&}�I�|���}Z�XG^hX�i���̺�a�P6|m���l(�J5��P�j'�W�欋e��+�K��onI=��;vቄ�}A�)�ׂ�_��]���u-�c��f��
f�ɢ���:f[�˱�F�(���C=�caoIp�@c�t:2�;JϘTC�d�m�Z�l�]w�/�&���f�8|ΐ��dD��{�޴���5:�.�w�ǜ#��.�ẍ́��\;t��3�	v~G�LL��דf)Z� �ޚ�o����i��D�E�S�`v�Ƃ��m ��9�3��!=9���~۵�vͿ``���ˠV�6Pm��b�`
�#l��_بf�OF	���3�H̚tf%ֺ��|��ٔ���r�<�ߜ�&���
k�
C_n���eD��'G�/��T�g�o�%�ʵ�dC�m1�Vk�Rm]Mh,���A��^�ҦൃЂ_ܜ��"9�拟���͕	�o#<(���@�`�:k9	��)��a~������>�+�5����(Un�J+���IĒ���m�'�����t�`������'���1�0I?������}[	�C���Ox�h-U���>�@D#.4'�'je��c1�7DQ���sO6!!��c#�h���Us���?��M�ٞ
(L���
(>�; g8�V�+�j������'_�3=CM�;�� ]f��@Q��T��N=B��?�@lu�P1����|����\N	���6fsoA/38��^h�:�s����Nߊ}���)�5=�&��0�*������y�)��(xs	1:�$[�����wp��9�D�����x��Y5!?c�;@E ڙe��`b0�%kXcJ���0�8A�Tl��뮼�^�skLc`�0W��-�� ��9F�LغVݳ��H��yn=a��\�ܳ��j��̱��=-��k�����zcLܷS5./v�2nlUg�m�l���ի�8� �c,��0Q�t��\9����Q���*��b^��5�T=��8nŌDʅ�Ͽ'��i�
��+�XM��ƃ�޵ �}c�-�}+��9F��읠��K!��W��lTҍh� ��+h��%�A�i44Kb4r�!��a�|�$r`�ua�b_|ܣ^L �'��O�K}�������V�|=��6�N!�=�s�xֽ{�آ�r�����#�,=��9�;������M(
�?��o�{�0VR��c�|����Ya�*�A��虼����(TO4��	��w��Z�3;�P�2��7~iIZ�'Bk\�\�H���������q�[��gto�0�*��Hf��������>��n�L��V|@/\7�&��j��|�
G�N�9��qY77� ���MB���2,gJxQ���߃q)~T��W�@/��J^�u�}�C�Bs�u^@A��!d�� �7�ˋ�gQ��vN=����q.jȣ�Ԭ�0o�r+�����Xv�D��{�@A���R*P9��-/To%6VmTK�z��r�-�h���_A�|�K�ݭ2�s�Рo�U����Դ3�v�}�~>�rui�%u"�|�7��*L!Њr\�y��q�h���B��rvqOĤ��u�BQ�;�D�TeǾ�/�
S�@2���&��VPN~_E�/�u:����@5冇l�m~�fͨ���hx<m�=z]D�k��SP�U�l��k��.1}&�W��!�[n?�٭�LX_92:���Q<��Ohd@=GMһس��&�
�cx��p��������%f�.��S-)��h�\���H���IR߱kdd�O�*>�v4*��	�ȼ؛����3��G�u�ڹ��9��#jA�}Z�y3
��9��ɭ����UD+h�g=��=$�P��M b��Ʈ@ĕ�+�a���c�;쯊��bs�3
�!��m�Od�ӏ���jhK�M���e�[��H� Sf�~��ZPH������i/��<�S�!�f��ٵ�Z(�J`��$7(Q��Z�r��_
�	NJ0�*�Z�N.`")��%бoٻ6 ���'�&[ ʻ��`d�1�|�@W{a�S�0Ħ�W	�����d�>*��0��H���Ԫi��Bw�o�2%�@���׵٠1�7��a~l��=�����כ5�ϭ�6�]C�*<7rkl,Q�'`�-_@6�%�ֵ;D��U����sv��b���$30���!2���v��@j���I��c��*{V��H�(�����.G^]MYv��n�g�T>nt� Ց+Utϵ�Ƨ��
���|@�qX7���ȢVX�����ݳ�.�tsk&��d����P���Z]ir���?zb�_`�#]M�g�(j�C�6:�=���#[� (���=��l���]��*۽h礥pa�+�0�;:	���a�A����%��s-���q3��A���~g���s[���1Z.���EiM��V�#q��bg`u:��#/�}:�z������~��3?�l��3
P]��J��Z�(\撆H�p�@�ipZ��7��(���2��Ѭ��E;�l�]�;�(e�|��������4�I���AK[����s��!v���{�q���M�L+�b�R��G�FT��������8,z�S~��N��;���Pwq���In5�^}�E#�����ЁG�>>|-T���菢m5b|�ކD�=_�%h�]�5���~�tͨ�Vm-�x��o-��2$D.����5^�ǥ&�:յ@r�~��{	���L�(���;���o$�����n��9-�V���W����D�
[����(>�ʵ�#ϟ'�� J�OWn'Ĭ �kj[o����m,�fdZ�W�Ǥ������E��:^#9  ����"G���l�^as�����N�I��NH�?ir��G[��/痊���1�?��e�WnkfI]���āCQ�B��0�{���}���_J��(���'0��ӥO9�}3·|H����+� 8 p���R��m���=I��m����e����; ]��w�<2E�]�k�E�l�Ji�:i��[L0���+����\�F����x�%�[���HE�o������O��~�����)N���]��rٕ?iV�VD�4kj ����I�%hq<-WO1�tI,\�/�txw�֥��/�d�gm��b*g�je�Q��zdz�W��$1_�0MRƀ�1��q'���Qn܁^���]��re�`���Y����!!���uƺ�]�$�6���"*�I"I@�~�)ӹT4�IN-d� l�})~_f�v�D���	O�SRd0N�ʚ�\����������)�eW���[�~ټƟ��T��+����]��Z�V�ʺ2��lw?�F;�u�j�ޞAs�_#�^�㶣�y�٥P�kSV�6���J��.xY�����K�����f������`iKwJ: �ǠE�ޣZ����*�#�����
��5GJO͵)�����1�@�vI �C�����p�e@���ʥPx�>/J�^鐍m��?�6I�`�E���Eq�1��RW@,챨$�Cu#��2�~5�S�rƅF��	�֭7-9䣱΋~��ނ-�j��!�
��Ӫ�Y�*���8LBeL�Ӑ���;^<=󃀝#dkc���|̳nZ	��eR$6P��Z��,y��� ���4hm|�X-�"�,���o�k�\�"ѩ��K똡]K��\��Nv�f?hK�TS��� Pկ��xD�pqAݤ��@>'|���Uc��);�M�.X�5�0���E2�� ����Z�9Wb�'�.m8ϓ,Q��]�P	�b�d/���/t��N�VW���� 4;ް� $~�vWHLp`�i�ڗ|	b̴^ts������5��pϷ|�L1���0eNl}r��(��[�os .[��U���bH4՝T��eZ����Z3Ӈ������� _o����A�p�{���7���y ��!����T�ןT:����*�Oe�+��ܛ/���0xn�:�i��q�g>s,���=iI�G�k覅2�2��eT5, o-�:9V���ͩ.[?5*D�d���$�&��Ea���x�9@�@�PT[���X�'���U�f���V9��g�R�	�-t���C���[X�v�@����GrA�w��"�0�^�Ӂ��?1�K��^�G��ʇ���~׮��Kez���@@�ΙÃ�|�:�*]�^�!�5CEu��p? � ��! �R�����/�JP��лEgV�h�:��.���z����(D'����p��B"~˷�G�Y�(��c/M��}�[d�Vxy[�Y�j���>�>�I~>+3�(��M�"(�c��"���*�</n��n'E1D�\H��x�<�-������^,���"�$T^��e0.7h��$�ޔ�BȄ��T��S�$���a:y����A��ed#�}M>���6�E��gF9�k�靐���T���*�I��[w��S���a�ʟ���p�� g��q��6ŏ��p3�� ��U��E�.ֈP��qC�=�u����G�?��L��S3�>�R��6�3obP��}H�)��)$8i]� we �9�V�Qi�tOӓc�ܳ���;&M��
0D��}vfe�~��ϐO����-�TM�ä�m��Q�����q@�Bj>��$��n�=����@�x�4Cgm��]h�S:��f��E����4ޖ~�+k�@�A;qv'��[�C���	���E6�NgT@]//�	�G��uвɚ�Zl�^L=H�B��ZT�K�N���+x[�)R��ʿf�\�vMBB�ha[��I=S8��uߑ�63^@�KPI��3_�ꆉz���|�Ĳ�ڢ����)�WK��	(��J'�VϡVQ�%�d1��m��l2J:@�RfeLç��]��[��
A��}Ԋ�v��Q���[��yC診��W�Gr�����隿l�_LR��(.����{�B����R|>� �]o�it��5¨�v�[7�.����&b� �ח5��p6�2j�W�y��&C���#�'yR��M�i��/"OݾZ�1�*�"���j��ʒQ�c�O��)�\Zǡ�}�\��'ל���g��X#�d�ʎ���v����4.�T�J��c�����Ά�;A���@�Ґ���������y�w��7�4Df�����x�Ɩ/Z�a����-+哦�;"@�~�-�+���g$tIڮv-xk�~�� �t�g�6ɿ��V����6�����C�ZIy�$D:�G�-ў�����fi�m�@4Q@��.頠�/�鮞7eV!(y�?5�i��'��^���LB��6݃������ޝ���Q�hH�w-;o��W��WoAgZ�ãfĊ��F.N��2U����c}�Sc�ϳ��������S����ꃰK鉜P������-"n��\b
�%3��@��x�ө�O����R��/�r�����B�5˔s^9�R+��	Uq�~t�c�0nG���LY��?A�����[���D�=�������:D6���xLs�n�\�����|Zni��e����=�~��՚�6X���n��X�G��q7r��X��E[K�JC�� ă؉��5�!ǚ�{���_�u�<�n�K�����qBt��SO�S��a(�c- �1n�pu�h��	߈갈�4o�Δ�� [��2H�[��~�<$��㥳��8������v�@����k��b�p�=:��J����G�ȋKCk	��
�|���%��9��;���}�e!sHy��'��BM7��R��J�сR�EB���4��6�Ѵg�@��B�H|�R���ǉ���'FY�ӡ@`�˽�H�׷wz�qP�Z���a�3^���0�������v�����]c�`���У��c���$�X�`0�1���2�V-��~l��;c�e+ʠu�d��G\U9]5�	:���п�;#@M�.l��?� g�D[VH]�;(�鮭���T���i��9J�.>0�a)n2�h�i|p���W�j�㊔�Zb{&ޮ��nf{��"�|m����/��1LT����x����/�qї�P��~Y�)��8j��0Ʊ4�>