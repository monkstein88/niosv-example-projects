// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
PGt+ejgXhtGmfrqCTGqmcxJOGWTT2iFb3HOR5gsNkbWyLR5oP85MveCUDDw37RvH9qQuF838M4DG
0KNTcJmXgNmhISnsG69VY4278A1i4dpl2RhnMi+sM/y6Ygt1I1bzOE0V84whG2rCavm+SA15esTm
tr2vAHVYbclJ5mbwYhLnvBzTO8vFCW1inj/yj5OUvXpcFCayAuhFBSQuOS+1Jgq2qEfa4S0nXNMd
EbzGdkY3s36/R+rtGbmFkOPiBbtmle/DcMSgse7DagW6QcLwfTo8xfo6zbV6a0FQ52fr7f7erF1p
/cviR/EQVGS46xd4JVJP0V9OfgdEi7MmMr3lfA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4928)
9CpbtZMWqnsW3+Q3nkGqbicgNH/r4hMxz/tq47rxhm1CigNqX2OjmAempDVQqRIEoL9nqKcuefZD
a0eUio6mJk8ZpSABlU/eJ+806SwoIis4+gsa+U6lsYGgaYWj3StzP8FKbIMJ+cEpryff+fTT2f4O
3EXGTJXwMcDNE3cmEPnAV/+vAu4JV+5Q5y1k5hltPOosb75J0sW8CcatCCG4jQURlie//Oli7hNX
nLU4k1WqzgUJnnO0LWP68wx78x21O9tC36CDXNhCHFtXfJ0dYYfnEsVgOByxVgPdMrndV2UydAag
1vrkenUAGAbyqv0tMOFjI8Chp9j6/YhKIXq5Uv/xI41fnQMMlMC3bP/Wwswp317lkzYemVTgCXEc
R5sOxyBIXPMGTaz0LIJHqGg7F/YWvPbB6ZODSHUHvFOJh3QaYH+EtGPO3HOIIns49sOls+WHSNEB
kdyfpN07gB9fsoD7Um/QOe0UaZsznS+/VOQVdTgan5p+Gbjk1tVbNGm9/lVqW9h6B0jiJhR/i9yQ
uNgKoPQVXLbh0QHykexkBjJCR6/LVeg+IV4FWJJeaR7tsaSTAAxfBb/E73G+ExV9GF6z3Kv71xTZ
22uvLFOKuSIlWl9V7S1ZJUos6B81K+QgCF2bfK+FotGFj64/T00VXHattOmfThM8dVRV9j9fQQpi
2WdsS0hRNYW1t/pkke9Cat//XfSuXq4Q2M1T2/I3FTXXPFnWKntcrZhANy72DH1WgdJwHEAzL0tD
BDxIu0bdB5fwV/Q3OpONkxkDGdqvYShz8vZo3nSN3kRtWZOvDrJuxJP7w3RdOZqYWkhGhUssQAXG
Wuzq3SM/n0DDgzy0K/0ZmWOM7O6bhchO7NjzDocBRx9kweFBfwvyJii+t6mqvWvOE8jqpAUoFCWJ
cw+BOEFfM74FBnZuSu+1R2oUUbGUrY44McfWtqmArQh4qs3mgs9DhdRo6sRxNPgU8JOSncwyd3SC
CS9u25UyX09SsYfKHn8zV0M2cOW4eAZ3zLNtWXgK7x6dTLr+mgl/RyoeCQohsmBOOd3PHKuGEPNF
U/RCWepRt4gdrPA5TC5MomNKHTMIub1FrlmrCjl1LQcXVFZFKu8qg4a57Fzx1rJBOnOxzof64pDW
YSao+HXjf896XKFuVMrYibo/JrH8qqWTvVSlnMRsxemWO2XeO6fPUjolJ/VjMAtx7v3xZKhQ/tjF
pi2f7uouoGQHqL60//TGZsCbIPfbSGlKP1L/Ryt0PV0L9sOiKcQIdzJuo45kk8NpYYl4/bkmXDlO
LCr1InZZo9/YGqHsktIR92I0Il9eYPzV3NddepjDpP/vh23kPJxAdQhV3WUUxIRPrcAn7otIMDRN
1uGSZV2X2ZUXMPySdf877ZlS4OFtDkcQ3jOAHETHzavqMn9dAOIhhlo/u8jXhiwQEBP+F0kR0ZJa
kzAoIGDh9L3Vq8Ar5NdfMY1pNWrKjbfemaoZYZ71dqOtciJxxiJK6srXDNmHlRO2S9RYql/g8X0R
4RntDDsgiWEmnWbW2jAPE5A25G1OfKExbUM6B919iv4weJ2tpCICdm66X7R53VvOWOrmexAgR0K6
E8mztR72czNT5DOH8HmFTt8/wfOZ/IuHVC4xykrmgYVPPMkA76bZzQZpyZJoOhHXfwaUvIi7Pa2L
VaZQ3RuAYF0U79vuIatzGbmEjDi6HsVyCg8K8AQGd7yELAG8dCXMZDnzcirH92Ar/WbdUlc3WHoL
lBqhB1bOkFPTnynmqqivdrwuQiCqVo+N4acNEqSNmbvXDTdVPvUGpBKr2PJm9O6Xtn9upZh5D5UE
BLMDeHj3Fic0ZxvaTNdIxsjdSqL8xiL/Tn7HYzpMxOKScLZHuhYw+cw+c2EUFCkJDAZJqnoDZN+i
OcZZPJBkdGc6JKx4k5WXw0j9vIIgFySKHrD1splE4WKN9Em9/CkizHeqES6foz6g8312eKB9wJC/
6in3AsBmw6ZmcQEGMmdjLAh9a+46klovQhrNeDdJxC+s4Utsy14LZWIbj3xgZts0FZYEeb6kGbkI
HECOltgcvFwfDU9S0pHo1IO2Nwa92KcqA3LECbzFpq5kiVJRnYCPjmB3q66B27wLbNVCdot+ZOsZ
oBMKSO7BRBoS2CuE3ZiV6uKG0r9Ergu8+K5ji63a2zHM93ZjhxHcfEYuRYfouY5hXCSBWG7CKDcc
OjNdNrBotahlwxz/pWx7cqze7yVC2KjG9WS63T0Liz54opYpm1KjRB33Q8XUQ9pAIA+k+6F9Xx9m
YbGsoiaAo2s7WCplb9ggtmW3oWl97TB+jr6qDHDiO5+AHkdRVn6XAcd4AcBH9Ctr58vs0877s5Gv
0/HFIr3v3aqyVH6b66BpiV4xRtrYVzOy5ZX7ocbgkkhLZ9OhEShG6v0YLjm/H3hxGGO4FzmGkARO
FL0gnJKohgW5iRcS126VC2IYm9URf8xnl+gCDWEi4weG9NfGdfHBVwrz0bJ5CVD5dFKA2/5zmiyV
To+Lym6TqyuNVe9GHVVI7HyMpL4ykP9v4GxJc4zjHsIWr/JaeIBrAUWkSB57kJL3jNRl8KuL/nZa
nBi+V6Asp79sxlEcomRbcbSU8hNqlnDwV8su892qlYJ412K8BykZCXGDmKIfRz+/UH3LcBoGTxkh
tl+U4BNjgL+gQt8b+SHqpnQo7sWUQoFEU1F3TZU1avvMVLNi6MF0egSP0TF9x0oD4zEgO0XIk/lp
ghxEwlP3OjRlXQwR8f2isySOcn7EIiNS6f5aL+C4JbkVSlajLWnx2aHYwRcmGrSNfJtT9w3B3UK6
UX6GdM8pEjFz/vhS91jR75YBeh6Ca4rB3c3OzehZewfwwolTZ2dN+Nr6t9OwL0O6gDZiXFq69d/I
qlAJzojxhJiV1zo0hR7IjEbZ7fjCIR2xgc38H/2DnAZz/mlXhhXLW5jyljRglOVyal6AHZ9mH8mA
j0/uoe9jx8bW1O1KIKnM0qvCvvaq2rHgKaFsdMQ1pMsG4MMGlurRLUK+ObXWrTP45KyziT5W9CrY
XHiTEFFGePbeG+SH/n0AtOPneYgkvtuPu38dz4p95yI8x/GFfaERNb0VnJMmkFt8VkyZG86o7MYT
f4gRyzmUrTge2+jHqkSU7dNIZPWT4jn/DaSb/ln2WFA+DtTuLVLUsxqo73EWREERxinNfMy1vo8N
ITPm4bRQ5XYFkHgWOo3Kr/Xo1mKwlZxpA51/CJwmwh8+ETS8pHi6AKySrf9PmjDrgoaupBp4mNHt
rZSoHGYNQUAyPZIm8ZlH275uLkOQpj9oEHCHSB7BYQChI4OSkcv9TCFpEzRvtxVZaHlAexxxCYwA
v+zVi30Hs+l5w7119GzUGdvv8CU9SFnC36zWP+N9IzR9FcUVNBxSF90TveYb9NeeUPwpU1u65nSH
yH5Dwhs+EyB4BqZfDyrEfz/UNBVi7RU2zFFyyxoa68zdSyEXGSkdQYAqlXWOIyRVaB2pnSw3X9K3
7dZrnm+4TsvQ4Ejn3CX+mNy2UpW/4ipL/JQFQnjEg96Kz2sqh1o4QZ1vqzu/HMnTOGPA6f+g9nAF
AbAjjT8ETMf+EQcrQvCO1vVhy1yDIg6zgwErjv5xpgr+kbvfQhlG6rb4OkRj30feRsu94IndAL+n
qbYSm7LhcFQU7eHiLXMh9UXhCqEp4tPBHZGKZ78KlWFeKj6CFkTkGm+aLj9+LelqO6SrkH9PaJMU
E1F4PZUKeijkwC/DrYVtUGbTZyTD51KipnQNWtoFk0sG1z/edoRc238oiYo83UbBUiDYwmhcJ+6F
Jy3/4se4buVY3rBzgU3jLUC5UIHUrW69Mjk+4Fnb61xaEvRkWADZcaIieGPGM3PsyJg0A4DevmMv
3tHR6ORwkXBIKr8QVpuiTmL+7ZtSKdP+ml2xPiQOD2TrF4udeCW+jWgK7icX7DNcY+Jr0coxSCRr
m4DaAVj94Gu3cK8XG3UFDlwLMjgyWlfbYen/ZrRE3IE4niSayvF23jFwGh04gnsE1slM68Zlfcni
dDHWWT9NJKBaLYGXkZFWHvfhiAfj+DouOYY8ca92+Tt45JCFj0X1D5MhoJsKfVpDpWz6yu5HRGXu
L3/iTRozzJIwHt4IpeTJKFDSrX7YYqQ+YTSVbwQtB7UCKFoYqDA6LYREK5Hxs7+2EpnpW17L5s1A
7I9GPAcH10QUXJhkM85NsE5ErhhfE/RRkelBLEKMFpEItwab8bezs0NwWryVl2GtVQWNjdvVUOQW
Wq6JA9c5kMc6Hmrp2LWRixrBDHT+Top/V5ePz1owxgQylLAH+7DoqxoVzAjciMMZlx9rBJFL9RN6
YGjDeo8/LQrH3vZJRenuB30aY2QaGaZj1QNd9GpA9PqxlHLaMbA6tWtO/T7FKXEehS2ghsy5TZgG
bJXmBb711vEkMvGRNJSE1+gGd435VYbqcy28R+ktsuxTzqIxIBe3Da9Y24gPWiTu/Pd3udu41egc
+/qyxdey2UVtDhzEDtxqGnNJ7a6/EDZ/UVasf2Z7NmzgpMtk6cXB228VzwIlVSc403bHVzN9MUlk
5lcMqtsqehRg3O++lNKtUsx8DDg0+9LqvqVXS13Sx7hUIlnfoCJIeQsXwDzG+Djm3wAago2qwTbu
KIg7zpufl2kcLWgEW9N1wm3IuddUKh6HAEya2T7sHrVkjPbWb8d6J6sHuXPrGVUFqil/bqWVIOp1
NirruMkj762qtIdGhYBARPMyj+5tEt6xhYQUitq5q84h19CKET12wULuOp9nI8KD/b0IzSmyUgMy
FCEBxDzVMgtfA8YyhZuWIAbR5KQhyxQu/KuR05cEvgaSekRHeDRDT3R8L0LZWx4BlQ4vwGE75Zyi
SZA3VbVrRYZbyvQX6BTJDMAt0vG0T5HFmrOIwEiHth9nK2OUrPAFkBrzjXekufdoAClcAhdtb7z2
VVYcEnMkLUHbpr4qDenu/W04Khu0lv3crYwWEBIb3ez4vDRVc+CQoX7MHWmrdUxMQT3s0qLBeEck
hxupCCBtA3/s664Tv5xSc5CLNE1AuKYWTA/Pllx6WRW5uV7ImL4MFi+C6j4N0niQbXKizlchvSVB
bS7WeNmGetyv/Ed68MxaHazGhbj4HaJ6OKRt8KZeQwXXy+qY7xuKbEM7dwszYitY6m2ljVphuiJe
D+FNmQNLXnz5VSoXJU4H1oix7fxy4H9iakPvizQ04cVij9Nlkm+UnlBaLQAs2J0CWfPm2QTiZfZJ
TPVYdOo5vynSjUJTTdNMXJ3RR4BHGON3O1Q1QP4XzKQqSuvleo2HEISHSg0baa9nC5Is0fbbTo1n
4/WV+22g5Rd9zBFRT31vCSTPwuEhXbkZqnuu15Yi1XIT6HP3wOS99Xdzzu4lqZaUHXduRe7zIvy1
1g9qP9agbaTd46NBD9/EabG46Nuft1WHrJRSGo/99SX6VzYhBlhIW2k1n8p+vVm/oufsPkDUOadi
rmQbCiLIcgL65jfrMI5Ut0+bHNM5HbC+gu910T1KNY+tiFLzOB6aR/37B6DRQEmwlPRbC9NGOlqT
keCYrOk5BqtZcO70/X4rwKWWAkD+QKd3vGAvP7iIaAoRJQ3rEuFpSVHVSoJNPgNNENp6cmD20K/y
Fz+eXsP7WZ1RnCMRya+rGB+HhTuYgT4h3IH/7mfSN3VqPnfxa8O6r/UJ7VSPejCiwe8X3I31gZIo
o4EyAgF2/AbpJMgehHzjw6+WHNCPDrWvmMkjPNvOSwbJz/N9/I5KKzboKesBY8do7JQ9GmHwXEUe
eTHzUGzdZkUIwjogeEMWmeOnxzlGS7omqJyPnbnI7O9WrfMP1CQbl9Q/vgddOi6i3ab2calcDB/k
5hBbNwea1TGLgQyKFyjpiWt/pOJcU5VxaZoGfRuTieG59Ud+ozxQn2z+uOEt919Xtj6zz3HGeR97
DY0A9cRtnTAjKRi7inD3EL4GD3UH6vcATtRo3qmI5hm8K6UL8G9/tTL+Q8Bb7igMkldExv2eknDZ
AU8aSMSfNrAHZcMAr89JOzwOrH2KyxLCWlgTUH78bp5ID9fmaD1fCBkTScjUlhy3MP14XrpzFVQb
aQZlme6jrWEQcJy1ywX2eeRZx79HCfC9BBxhvRRqc6CGoHBG2NfDB4F+CKbFk8495UZW96MTA/h/
VTo0PZiCsA/M8pJqbtrT/JocqzhUF2Ygl+SjMvoCNGgoM5bha95GIL3L+1tdmlnI0kzigcdYjzYL
de3vwRRJGmm3l5Jm0AAxm7cCgM/F4Xvt9oT15kmUt3i2rcaEC0eFKjkunPV1E8/yIS7uBN3VdxO/
bDAYJ9WZ+tsUV7/kSqOH3DHp1MftDecJFQU1lIsO9oodKggvjBbvoTKkM+0+ssbKF0ljHWvNuFDP
pBsP3haAbHjmxB7o0ANfTcamdGzB7rdMf8JHcPjvh9NDwRwNAkyYUdKLju7uRLxoj1iDGXp5NL+g
ybkyiUnabsmpvX0/6VtAaRS+d8iwA99/5OZfMtjGI8LDY1SvkokCzuXs0e/v313fU5BcxjAff9z9
SBUOjs8GZnc6AfHXdkL4JGskkHDV9qfEGUI=
`pragma protect end_protected
