// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
m+zWzHHVCJnaxJtaPfE0bPJgdpJEnW6wOxT/1BZ1NHzWm8KxY59zBnJSGhrJ2iT/8z960/Q+q5Qe
OA7gjk8p+2ZErMZSao/zukELjTm/N5og+H9QOFuJCSrT9RMn+LBGUMVtR0txrume+c+JoA4fnCKd
WoJNEjnzR4zCKFtbSHT20g8vtTeMchR/w3vjcIHo24jZ30ZVIrEwj8DmjUxgVL4Ot04F9khncV/J
C5Ma0RjSjhq41YurToG1APu9utDZ0MBsXSDbKuK+PzDKcmmBpO+Ax3lGOSXje1IjBCjLN6k4WWhp
ouFuz+GhheU1zBYIJkC/HJnRP6jNEu49WGDNDQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 48224)
eHZip6MmRPvGw46tk10BUIuwFACVI+YN7j2T0WQEslhRC3YWPYSVY2A1aBw7E1h54peS+yOcki7j
wujxeYpznijb4pBWJu8WDFFjas13fKJ/iQowlL1/KHGpg8JL/nbLf2kp1wiartU8435eBR3HgNGs
dIrsmIdLl1Gsky1A2bL2XeaV4xS7mBCkIt40VCPvThhwvnPTjyQjw6cAyw3f2skcLqH5TfyrqH7u
j6jolWWz5MURb82cSwX90wEWYNdv7E6y9GG5hBSwqgscNDkch8kwQUhTxBq5kFhhCnTH8UMrLN4P
QxrVmi7SW6YXwdgOrhY3QNTeW1o6881qS7qGENpHzdBR+NNTLGhurLHnmw2uTRNkE6BBR6PGak9Q
mx0UBJJOJ2zdPD6fzveYxLg4as0ZEJ9Vl+w5Sj8GBCuBgWTKUD3RUovyXA1PFTgNy7hN3e1sZ9Np
AIm//y0E70ccTbUZ/colOKngu9kGENq45+uL5ZGJgbZFsbSuTV1F0XF3ig1WU7+OBTx4z5TSozPv
9aHc8lKSrzR5QxO7xjJXHxw+t+IkTWLpjI9i87K/7dXgHehrXFosisag5wX69/NIjfVsSGYYbi5Y
3/B4Cg2ulidPIqd0OtOsnbb4B5oaNwnMHPEd39fwcbeggedsVE2bZdVu4fJtWvcgJ34WIV0hWD+Q
ZsgQJV7UJN4Z7P2pUr3uv6NUgH5O56GfZMJp+tl53fa2Pj5U8D4Jthj5ag2gLQTvQXXvVSU1wPe1
m34gEzZMK9GwDX3Mso3RIvNuUYA8CrWRx1zafjcVR5CnZV1BodAP5YRUaOIE1/5yQbvYBTjOjtOj
k5g6+UCS5ntcResm2fhE/0Ky3cM5YgkvEaL8Avy06HzLyVOiMlT4ZUQTvC6AKoSHsgDOoDzmR3hk
b8OWDzLX/H02+ykMNKX6SQwKzP/vWeSyhFFU6kMO/bwNIX1EHTyaQVrP55nibCOlCswt/VcCdVwZ
2OuIt9f8bLpVODhRuo+4fDkdOL2frg4xz8M8cfDbqfvP0QcZrGVE3AjjNGPu1ufn00fwiBj7fijn
IJ/15K1nJBxG5UK+liwLBVsiZ/1as45cPG3u1qLFoeK6oEmIIf/BsfF35z7KfpPEisboofROkTrQ
tbfN2BptYxU1JAhKMQmP9OnPLncw1TGdQ+aT6z4lBQCvun/++OTHhYhZbLq1pglKUm+gWWsJQyr4
vz1bzoqaTTtN5DqjgvgwbGV6t4ZOcR1LYUAj0Eo23g5l2v+2XpHI1Hbq8j3/CrPaWVB/H1eCqVw5
nWMYGKZbfGve0l5L9oxJn9ADs3UWoDOFcJGzmSASC4he9JYlsiM8ttC2OKldf1ptJHmVc5lk/Zll
v+UDwApxSRjnUpGAZrfbIFwS2fpt5fwmm3IbGpbQcPGZxWmLDegbtBhrAwngE91gBeOQ2j/4e4pj
6LFk1xhW6+hByHORZr0oqCFyeHbA0DKF94ZTEUsZGvvVbOHoF3gkz28sBkPJ5K9KnXeXfJd0xPPz
SJnUZ29mp4FcAH+rhXx4y3q4ZP6BzrlI2Mt2Ca+/1jbM9SG/04WDZg6pFUUNgb1SBftRBbtkLQ3A
dm885PZUrUf6cCrQdFoMMFZLfmMTgQOLv2qobUnxTjSlHHmu+fsZ0FNEjf/n2UfMzgeLxZHaymra
YCzfN3yFAVHVGVTy8fgznnlv+g3UHrA8aHfVNQk6m/tuRPToOiS7dmbjQB4Pu9ZpgEZMtmAD7QOE
yDucNWiTIyPNiiTf9/4r3HR59IOR5Dusf/MgUlXKD7jNOebMcAy2zAo+kdWg6eRcJzBiyV49BkeJ
8L5WeETGai+/FQe6yjBAL/iVqdo2Nzpm/DQf5YpDuqIoLTSPFfpJ7/HLNpnLi68F6aE8MtxcZUfI
HyyWps/QPshJpF1yXDJ/bCndDgDjTZ37D3Fh6hYWUItPc0opVNFxp0S9ev3FRpIS0yGpj0M27aWk
kgntsmBM5OzBh7NkdEXfkkqleGeHRoquH95RNVaXtrAwwlyETJ1b8m8KKXAptq0PYkmjnIKXUMdD
Bdq9khF/2/KU38DRP1CsvDa6vM8jwhfePzA0AwQcki8lcuYqf9hf4+iDeJzJOXiwticnCvX8G9Ha
1SIO5v/ao9Utj/Jsz87kRRQVrZ4gdiPl98NXlFiVsXTwkGgtgVa7SMc6kslQCI019MS6B2SBRhij
O9e67H6IE/7y2N0Isrb+ZSqZ2D8hbo6+8bNzq3fgzkwVB8QPBSDvvsf5kuzrGKwKvFtMQoirhl3u
gN+n5yFxBsnjik3fb3da73n8RdxQCSO7bY9yS3dV/gXtN/dMtqialISNbky+nCZr5NKQYFhj8u9n
gkWEHOKzlnfpYK3HyhKzqGQjEszFjxtscFmAowc/e9byaeGpAQTyc3hAjnuhZjbxnH9QHN5ZW3Pw
DdHqgTIXjHRdHK6HkneYvQUXHROFYPpsvQdGrbcZIWrxKQAoQyWPxHxfSMjWGLOECLeQD2Hm5sZi
5rW6PZtu4Wbgt+RBI9zWMYRp07kLjXW4PTTwbK9PP9UTj6R0nOtyb/4h8jEmJl504ZNyHI+UQuiq
M9mT7QNbLtV3sHQM1ZO8+3D6S1Ifos2DCljfZI0V8Nnymmr6xXTI+RciIFrfqQrhSlFYg4PwCUwq
N6reVPBlhaVuYGaJYeJClYqlM1mMZLyKY/gfn4I2pRZJO57A/Sr6zeSFRzsMH/XEK6OZNNK3ipWZ
/65fIZ10MW9md0Uyscv0nTBOE6TFJUFbQecKbVo9BSRf9XbW1xa95Gpm+woGABO47lCMsDQAqcck
m4jVUAurxhdMT1fot+468tYkLy1nt27AIlaTe2QWCFBivIRq/9iMCE1MH9TMWeULOPfxVadR50Mj
oTKJuz95nBCmjbP3FU0wqXlPGloE1MOyFlCDNe1rNZVCOTnx1Ly78hh5aINCxMX6K3E9Qp4JFyIX
SuCYIrckd6N9dLJCk5U8xDZkMk0Y1HKzlqSVcnNkmr41a2d7gW7MFZoK87SM/ZSdBqOFZRFk7SWM
LvwEkyLsFhR99hTXOLeZNDKt7OeRHOuulnLS1YkUY0U8CAB0JKJ1QDrtIAd0/AX/elf4p7VeKURL
GWblZeEk7tRvwMrHFsqTCmdFC8SJmsQRJ35hFS0I5TgiJr0is5566AD/usC7tCW7GcFRitHSj5bD
N1Ljk8s5XRJ3uV9Ca77XMkWsHo3irZDJFjO0IxwJffol6hEVzdpHuOTr/sJ+aTrYx8mSOXvhgH2V
sqltOJhNb9vS1TaldPCVYEudYS23dWC7thXUgRtxSmJtvui6S2nl9Nz6OcT8RGpmp8WVvY4xRNo6
ZYdxbDs0dEbSWHUxAfMwyl5pqsSSrQDHxmZYa7bjDR957xMflYA8u/SGVxZTVhu4zOxpQdD2aUvz
29ggrQ48/khn32IbjJVlaJ1zHME1pX+DDfXnHYKRFghd/CQ9VVlKkUfc0nPAe13/RCitk7KCkewz
TI8LxPDXT7KG8hbvaHTYJtS2Vek++k0swi0Rx3D8x5mv/rEIuuPWYa1WH78vStK1CegCqx6GjmnN
ltDRmQcMzgxitlq5iHvTmhXbUkSmy07+3/FMVzHX9HREp7L9gD96fHuQT7XpPZPi0u8CvktM1Z7N
VizS+ehhjugq8RGQVdJsaa2b/E9HdulQnI/7EvZ3y2wRah9XVVVe7Nj1jHhM0dSIUjX7E+QSbJSi
L71S75mDb8l01AhtzSh5LRLGx+rkanHZsyEUZee/dWMFyct8ZBpgzLRu8ojoyAuVRwmNUAHWa3g2
pQUK4C50Fftm9NDzpzqgiGCv4Lf9NFH38HVoVp/lvLLBjkH7ttbwl3oJIRP10Xzy11OhgtjdJH3T
HeKjdvclLdpNxr+t44ckOY60YWAJDSGP8NwpFseIifCGmnaUwMETXStaupVRnANVGA1h0qx7DYVE
UHeANAoh9VmOhzzJOqGbNgN7V2Zk9DkzOVSrdH4HPGD0uUxTQLx9BYrHd64bjS2+sWIuKJ3aTtoR
LG7yRRH/wDnimGjv2D6BoGR/UEumrEQLsrW/ZtcI0cy7MKvU5XlRlzx1Mrh6I3JCBZxokEWNBWt5
afG1RGnccvOFY0Mu2uXoPpuMiHCpvfCfVu+5xwx1MVeOCs13Omfw7tEVWJltJ7z/tOVxDM2xuvRQ
UXskIgy4wXb+GpE/3AWogDJQacIBjnBZ5RAGft2GH4cAQNAK5QC03dx92TPfgURYVCxUQMFzn9hn
Fxc3YmoPlxNH+3Px2aYZ9Ezr4f+P68WHPU9Y/w44UYSLQzcuZmfq2Qa0eWxJtx0gC5CxMpSenbmu
qZ7iqomgqKgWrBValc4XMj/pvyK8on3OeWYUEZVz5NYYwUoOf6vrp+oSEvWL+KJmvU9YgImQ2kiH
kMZtkF+jDTdDWO4JUl4sXmOC6ttMXmjOtZSVkz3KFJX+WpZBNC9qdkTrBfdhschixT+bPnIXMoIS
IHePlptza+PV5f3SgpxthJjdE3nj+to4da250a5y1T/9cA9YVFky4lR18aIcBNbLh23AefpqY16b
xQKt+RHpnQqA3IRcuu44JO++miEJkcn8hOu39gFFl7hQb/F2O/ODh5e4JPbrKQqxIK8YmoOv6i9v
f69Bh/+R5KDf8gdad6aCUmcQQB5Z9HQImWAJ9LncgSVnLtiB/DggKFMXVgVYG/40Atsm/yBcs7Wg
+YiFhfztSMZH8UxuKGRCorItU0ovZFVPgE4W/vzOWw3IqmV1i0EW8hdDyWRMYMygr+GapqvsPcRW
1s2zzIlADADPNnsLfQG3vffz8/+FyPOwk+9NVTssjcZfTwrq+tG5yYpGyqDNKnUdsFHN+3RCVeDa
c/mcK56/BZUS7L68iTxh87wshk9My0Ff1rQaJd7CmKEXY4o3QUnnFWRfI+KvRAkUY+1B7o6oBYow
UilPZpMEShvfKITlO+8cc4YtIS4/rJR40PQak7n4vmT1TnbRLsZ44XCUWfhE0FyHsrfclYnaOjeX
/YGeENVmQDEC2oZD/EuHPgQfSFCWsu0xFxFKRqMjew6AtRp2ssLzUpA+XKY4FU6q6ZPZSfvkrNL0
DOVc04aotNdXa/CCd+QeDkeQBssRBSlHkLv4vl0HLok61aHHnIUczSTndFgmoM+f+Ggfwgp8tFhV
kxYfamLrpmbLyToMlmB0ayvAv/wha/NMaSN8KygSvKOLKUEsyHp4rS806wYdDIrNs/RNJQKfYHF0
aYKu/c/dkA+Rg89geh0gPmt7ZaAOGH1KcmxR6edoG8YkKoN3ZupqQ+ShjiNP9T6KQc5EFS9OvB4r
syA/YdHFzOESGS/XUtRFIWb/WeumLCiEJmQRE0jLV9Nj1RepT/RokwUHfy7WR+SAbj55iFdEvJ13
99abvXESal8PSl7MInyeIVwTMbL1MJCWu5weov7dEBiRBwxZva1s/zi/SzwZeMTpWB5esKRfNkuZ
IVADjKAnLsYXxsT5hk4uzPYW54EQOvJRXahiL/oerrVSo6VeXHj+KjsieWgcvVoqLdnjDMQWW2eE
qId8PgCVZS5bPpkn4sfHHfBj8e2LYAovMlYkW9Gp4mjfWRKf3RzB3PE3VbGAOCAeJ6JkKo9fij3q
6ArzksWSxfi3/agdLB99IGwFVgQM9NH14PmeiSeKbnqwXpONNnTUpvXPf6xvHvkeKjxzyLM3MJzJ
OwpEI7aUVTUcPAING15vW5jJTYnzmdcLJEDyF3YQT+YGeTHhYlT26SdhRALaU1Ne0HeF9rd9koFo
b6BCcn4CXLNibXbnY+tRPDhPTy7Legj/PZn4L09Nats3Rjd7Dld16HNqkes91hEN5hod1RIMwGp+
un9bGD01UvCrTIGfLNBVqn3uzCfvKnOzPzncw3D3O1XBTp3iDTSh3Gy6yzxkI1uqPljfAUPqQn4Q
wrrPIydrZyDwRurUetYFU90upps3QEFyMGZV7bQ0Q4uJUmDlZ8XLAlM+2WKwV2A2sSyCEaXEvAqt
HmD4jWqKtWrbwXlztKUxrqdGd4CPhWnkuKx5MXHnGGwdR+MGVho8YLs8ntzayhXy9HuKNGxIXGUZ
P6ldlHUbDIyBx1PeFHcTlTnW7Rf70+Rum6laBqIbH3la+n3MDYAXNv3OfchmOXj0cAcEjJteJNJp
HxovN50TDNra6sP/thw1Az8lUAalw3pS143L8Ovp+AqcNaXI3sL0Ziak0K64xH3Cii9Fb/t/YWIy
MHnGoYzmFvj6V62RAkcwmBeX0Ho8yDACNozLysth6pNQL1jkCS7UjJkFu41xL16+kLEYE/Y1thJ2
z/KRjEJLH36kCAUQ/TqGWEcBfeVntu3SMdY8Vl3sv4faPJERe9YNweGgkaXkqqTARZp6SUGhh33T
nYi5ZHUJnewNFmiOLK64YxIWrqX/SxUd1Pf1TRNq/9Y/tIilzwZjqVSlcXXEPJaUM6Pf3cCgUB0G
yuE2edQtVom0f1uGEy3NvynNJKjk2UrOsCIZjz1l6GQg4vg3s1Ml6zrK6cggBTdbD0Ums3f0j5eL
HLsI5XhD/FQRbNqv0jAlfsliV2r7ZrVwO1fBKih76Njf5q913PWsBVBBZEeKUAFYSdsvsTOCIKB1
u7pUGUOv5LjxzlmEiUa1pVKlzO7XEiDi1nMKWlu2fujDxRQPwTopEJ4LWqIMUP4Z5SQVJ4hc6Mro
l9pLsmCV9vicjbflbOPeNMALnk4Bn95Onal8EZcLr0VidrHiGNSDCf4nT1MFDpnib0WryQ0w2AZY
7CnnvU+n++Fw20F0NZuqXhrP9GgtGG8qvoHgJ98eIaNaVr32ULwcxyqt0i0YVoF6bwYP8GTRThNS
wQfdjETh7gQsMNPzUbyrmj8oyd1HfjfGA4LwK98mp+oI3ktT/vKSYAU/54T8084SV3NS5YGk0j5R
N5YfP3oubKl0363Uc07FPPg1IxTK/JMaPau3PBKuodP7X04KrqK/JxA0ADcnr75S55nX9Y2F62h/
nRtqWmmseT+6nhNt4dTjZqMJnAY+Luetm23m1cOff6zEyRinEg7GWzaqE2bbCRQKOILn5U8IFRJJ
LcSDevJcNMH/K70nTozJa2dfAWSLi7Bwog+xaeBBFz7igXi9LVFYifNhMahfTPUSQ+cjII17tgk/
x24+iuilz0mvO1BRYCKC7vDps8Mk29B9EASmxVXqzVhy+JTJF4TeE/8bvLV+d7+UE21T/LmbkE+D
cfN2+839PHk1RgY50V+6tF4bA3vrKCGT+X5S8nGvxiDbDTNbYms/GnHOb+TVrNAV7EmdH7qyuLZ5
TglcFOVAIgN9BexPp3a5UnVVMrHGJDoY7wAMMHjGHwtp6MRRyt9OZoFv6/QC9Ck1VYwlMHOFmH03
qFt8YBktGBXmIw5D6KxJkvIl+40eIvobtWsPROw4SNQCy6mHETT5lMBoEXh4Kn5YW43Tc0dtp0Iu
XLmLvCETE+dGOsxRSmYJCEP5Bdafbxd98FZO6Xjadx1PX07WMbsfzoAINy6CbfXe72/jC3V1PJ8V
chw9P3leqVhOVytuHim3yTwd/EpLcdlEhdnbWOezqxVsndMrjGfr8lwTonRY8QS0/g3TpBJHT261
sNNJZ7ExqPuQStK2Np3ArfwlLfVULxWg9SWRF0ye9oqACosESZcq/1MBEhag1gszookQijt0ECJY
7CjYm4dOOTSsE/phWhTTpoTqdhT1C7VmDz3TkbgwOlkZgxoGGFdcamYD2T5Xk48EpclxVEUs7kOY
zwre2dbb9AU1KFXA2h2s3PzyP4r0DsTWxYg9Wb9YLmDIqBz95Xs5XhgmVpaqxfigRmMCPTRucXMT
AZgNgCOjYCUDGvgbKaWqlihlWjFwBxauG9eSH0UapWPlB15s67cbZo3pJST/PiE4yNJrTvwSOpOD
HiiJwk+DVTkjSbhm4tHIycuuCXHfiFuMyaLeR+ndt0U1/E9vlefIhKXGU1XZSs1kcqiR3mlwJwhO
ldkawZnbmlL82DYqLYfaFw9xDNJHRPA2/xBFg04RLkwL5NNtEy5vdeRpqJZTO524W8TcedpT0LYn
c4jahct7Ktdn2EugZESYoqow+aKDKmxAtZGenfw2bArPz1hpVLjWZJfus8CHJNHqKqK+dBw+kzZr
dWOrl8LhJnp4iEslDU/DCNBo/3hlhm/M7pxlaUjISlDrqvA1BGQEZT8g4/ToIzm+VPrS52hJjt2n
NVq5uPEOhgxS+KXyRnBJXvmWF1amOHey60fVi9KjTOv7xLgg90otZ+3rojCJJoib9TK+6uO5Xi+T
DHUNNVJjl/br/+51e4Wj9eihLxWpZCODPdZdwJ+FPRYnx1cY1mCb28y3BfAJzoKKlCllyhksU5OM
8hpBTxbnqnCoiLk60y0rRWKK6bqujgVpEz90VZm5OLKbEYAYPQeqeyqVQsX2b9OBHXQr9LgMwwKA
ztqVxb4G+ikhkBAI4wOB6aYb2eAGnaFuBgGUm5uaiZiQquOiMoKhVmi0uguRp86N5xilOlCAvrB/
d2YMYPUYHXpFgV+BX2btlYzP+iZZnDjiPcYLqnGjjKs4QczrgUEVvLcQPtWVxmObgkZyKEuzJePS
Lx/LN3fO9PX+gUcGNCkmsEz2Im2YjknnUs54ESL8j6nBjq0/JQb2v5aZbL8evnmksi+I0Md7fviM
dAYmAn1g66hi+p+JLigbiPTtcCFtZ/DD/GOubeU60EQ4Z5sp07ns4o7graGrIBaUnSD/S9tYBDEN
ddHAGQmG0a4568P3B8zXdTZZlwPT7JM4Mg96L9WaShLgmscGGYDPo0xYKomWmsIohjeCk54FrlGb
6FVABpLU0Fv/ZNCdxCrzUgAXenKf5pp/3vdWDuzh2gBwyRazoBN/AWPFG+Lc/RhTWtaBQK+DXjhV
q57lkPLZBasSqNPTdg3U/B/929c4Nj42LbNxuZZN946K9FoKPr9kWs4grF8wodMSH/TRBoIPELgE
8OaeTE22I1OgD2yYYjuegkHgXHCxOjaJ4QiKEzVoPRk6nK67iALKbwFnEpgt9UnDD/T3MdvGxQhq
VKYTE3t4oMB+OxgoiszSr/Hi6Ud2+6Z3eeWNe9XkkVmwCEsXmaOZqUpsz5FujcDhLYjm+eEAzGsm
R70qjjsqVaD7tbsypWNtIrSGUmRnqhAgCTqJd5wOwoFK1Ej6ZHE7lbfWWZiawjI7VY60PR/L7++t
Swwk7fd268in4EPO3yPeZaLAT+0AksLLF7JDz/j5YyFCdfylsBThmtVqvaKcpVGdRzqRgNyyTCNa
H4HwFzh6bL61Y9Wir7IIS9xvSFHx5CtqDexcdoszfg942/feXU/04HKtK/vyhktbwfi85lI26gOO
0GeiftjOA93aOgxuC+CczYVSNvmjPYclktfliU0ZlBbaO8ZYIDvN8q8d/RcxXexWzv1MOjWp9IKr
CN7ciyPD3+K2Ho1BnMHS4LBg4P9TbFxorDXzpLo+/5h96e1u6sqMFHAbl1OANsqszCMSuyLx/gR/
nkP20L6bBqFE2KMgk35xZm78YcaPT6p6rQ96w3GD1LFNpktGA7PPMGzuWY4WlDhNtvs1LsD4v4Le
tHWPX0x0m+9FDYejDzdiAIqK8sCbm8PeBsjLB5zRdQgKUVVboIw2rqtbmZltWmbwOcQR51HIcMT/
QONhF8X3xVyYt8mIpFee0P0g9MLK400361tL2DcT4hnJGdCa5Su/byki2xTGqHUnzzkNFRPQrxLK
QL2AQo18EXgi0dNUlDvmYYaHaKfmczykRSFFouzM0NiheDV3VwkjjynyarUmk4oZ+GJWEyjfjWpm
z+tLinfF1eTO9JVUBS8jIaTwmU9GYwOIxWYKDe5lSjHhsdRWD7haJDbe5OOIPxTZazPNldFR8BSL
1Q7rifIThW4eSor+T4On4kIK4hRouELGP4c/lvB8wDql7uUBFfekdxspHK4sZUxLwVeWNR1Fasr/
gDqtY3yKP8HI8OE1IMbF7cBXNBN4zbiV3uIyQYubrAFYwxRRKlbOlpLCB2nYKH1kL3TVO5CdDz7z
5CpQ8l7MhX+Gb8mmhP+8NaVQPDahSC/hXrSlnS48zRnZPofZjQzRPrIa/32MKQvwDAlNTO80LvvN
jEC1GfFDRm0W7bzUWaZs5CQynW6uC+dHzeqp2fNOOesyKkJjmV9Z3lz6hPqIXuPASQbFshU2Z0WF
WVHFdNRJb1zTDptZfwsbI6vVsV67WBO70I+c8aum8m7vgjanjl2C2a33+IkKoQhiunDO7ALjr+RV
C4aie0F6Q0FXhNf9d5KMWc9Y/XD6rnPFKVv0PTg4FBrRkwz6nkqmWEQTceQGBq0OfY1MfW5sqHLG
i2zcuVtNmYCljT0WrrA9uEbq2MngK+VCbfNjfeINq4FvwmHBgUrG+jCoeZLBf08MAD8lqlGOQuxW
AzgNVMKwAbZQawf9J4sxP9CE8mFtWzgCD1gSLUjcvzwAF6Nfty0y9LmV5BlBLNcRmiGjo1iFb1E4
dJ1+NOhsUBsqwghGhraJJeUSzGs6MkBMvNdtLP6wkQ63fV4h+mHSH3fhPUXZS3nVSXUkH8N4OUU9
kWFvx8WgaM8bkT4VqSvuiaICRnEtVFI8kKFiQVamg/4UpbeUEWMoakhieDW2WOaU2ddIfqDJ2X1G
i1X43K6tmJTRNq6wrsGfvNQ3h+j08a+ab8RT7EGwWFgyR4xzDPWugJSY3XA0T1PcFcRBeDr88/ER
LbeRFKZaTiv0OWCjcJLiMChZCyEzfv1LT1PGJsF9KGD0WMy5WVYOvb0tTLVm4f7+ye9oWS9f6KfF
oJtHn0g9gfU4CzqehK2hgsU8snL8Wfg/mViFvWNTtIgDTgXsSDcxEAY06Rqycv188yLQBJdKM5Vi
oPX1Yghhghrnnqx3YchFpSOpgg4XCtDWhesX+t0ytNgnog3aRqWb9K0fMhZHXzRmdMYgufF6vOwj
oqax+1Ma+uj11mPTqccbDi+jlQy/DKavRSyNW3WTOBs8CPLYHGj1/cZi26PqAg0xyFE9/s8BP5X3
GXfaIuvmM5PLIKsOyDA0iKr4JN9ctqB+hYhOUX0e4/VxqN1VT1rh2iC6j/ur60Ud5MFgdhBxxTrc
9+Ss4B72h2QZGsAf4AI7IkGDsJoRfv0J3dPv4K8u8T0sfpRDYvSIFxWFeD8QFeOmmRoUrr2FbqKy
atxqjtl8nmM94pOmgrVcR6G5jYBgktnbRulQsrz6hMHodApMuAYxriTnEcHR2CTlsqX+QEBGnyUe
vS1bAFs7VHwjMC8dxfQ/PD6dJkQE09U544M8AhyPUfOA1c9bv5FpG7OMyZO4oKjxqYbgx7nLTxpG
I6WyX0I7AQWwclLYqEUfDKSYsZpJDfnPMvCKMGeJy9jRNw0d3ZInX0y8r/ltOH7Gr2mKmvh6DTuU
XFczEknY5mxWsWFAtDOYxtbo6HQGvO7mOyUiC/22fXRdfoUWjK0YU8fkIJ8YrWkrkkIAAhSXQqMH
ki8Vzhp8sC71E0XA0TTyK8neCOGTilLSi9vYuOSOMPK9wY0/bV7tAPkBAN9MSI1pZrLiYUxUf+z5
Zjer5Ss0Agpgh36ZsjaajxX1DCgmyk3lbSUfuUz0QYBh1uFhMmsVkZTXChjaUFwO+K+5jXr6NelD
Vf7yUbad1ZoImDr3OanKzF84mwQb3mOqyMQ+QJX1M5nzgJazsrYgV4ySiYfBjlsHLsfJ3Dyg8vuB
caxqP3Vq6jkHz0aJbDdriwfu2C8/k+UX0kFnz9uYUS/Rqxp4w9q2IWdF/isCZpsURHp/aCBP2AQe
MWaKLxYW140J4IwGiJvmMSV3QojRABGechzHiXUthZxteTVLo3JrXDcfesLusCI4Q8ta0SVLt4Pq
XR/XRDOelSi5IJxjaz0cW3mPa2YmOewVyEd8GwAjMlwXoTXDa3xaON3U+6fgiEz9R4Ps7s3S5sEc
j086Xdcpa1n1rgshRnEfZvubHcwbT4f6C1sTkIf/ReEjCiB10kjObOocT2dWEX12nUOrAmRvTN35
yvNXeS9ult1uLr/DndkaMWVrfs838IMQxHFrw2b6zHJz8kdeXh4wH9zYQjNtIRmQk1VkiRvls51m
XmxWWSLDwmzctNJa1gSdIbnFhzQlkV7C4i9NDY+FXLh49mbQawfqzaZIjbELNW8R9oV/Vi8f7lSi
Dgxkp3Wr9BPWZNI7ik/6gBJIrv9qOO7jA4pljrhfe+MEHTyVC/c7nqS9U2fuvR2mLtSLqx9a0Axr
ASGb8A5Lzyapkslh9ulsHs9+uuIqc3P0MzjjAdWTeVcS49PQu6ZSemHYij2VtE8jkriQ0RNAPmwR
/NPG8Cka1bOTq3EmB3buGvJUpvLBX9HNVsderRSeUSh7vBtKcSsLcNXD0GJZIWdWSR7FqHelTSFA
S67DOiZGZ7+RV40sNZ0VlrVKmaqiLK3ZTZr7j9MLMYHYXGT3UPIckhHs/KBEkbg13frpyZqBB1wm
fns1RqHhTXG5GxcKvMcxJu09ijLX6zfEHNdEBZioAfrCBI7UcXUUTFQtxRYsHxTGA7sm3ITm1YZR
pIXyLV3Pca49trOpWa7hLj1nvHaqlIqKSczWnJ9rediKkn1w15QvXv9AelbHOaGwsVBqLhqRECP1
P761VCKL+w5DliB5AS477+1aBW/+444g+bAL6v+g5MSyB15u0CTgBNNWzzRQQzZUNV9q+Uvpkp7S
ZIW40crnSfOGqBNOHJZlF+ytgIjcPdE4vNmJ5uskqqE5PCV4nS9Gv+wyNh0h4IUlwl10g3NVYlrD
afaYFXZXW2Is149u8IHa0ISk1/+MTsquy6kLWorBqrC7cB9a4D1HqAccEI5CPNy4tQTDK+tnwPb5
4LpfjQD+YoOnbDsgC0pS2EWU1w4jx+93ssYJDJjYqxED6YxPj72vq+Kp3kntAqwvICWXGcqNzIu1
teVEUPEqU5MPuwC1/Srmpw7rwgOlITgHZrZXqiZMKRiVGlpZpEdZrn/kk26Pe6jA8ohGvSa0P1GA
NFQ6vzXdaeMXiyWCjIdI/2QV9EDyUXgm3bN1Ev1GCnzSPwJ0br/XgNBnCIXMUGNwxCxdJ9pqPbz/
binLIS6cj6aq8O16d+aNziFpolkS274APTymjhQIuhJpf0pF7vX+YBmGQXH3fz+vBCNE25TLPGs1
TELtcKYD4FPTZSw/vE0OL0bLVdXKdXNlyo+J0wR7wIS9wytg0lbLgVJ2JzeX2A6mpQvxhSL7zWz3
6RGVvNbBjDB8/dYLVkvEe2mf6tarREP2Mh6uSVvaA/EKHfmB6NjCtPzMrYZQQzVi9RdVCmrEl6Je
G3500L7bKtOQ31dNJOa/bKb3/x/Kl7kAMpeCuxfM4SuWmU8q1jyEunYMKIW3eNUjtI3GINNJdkp8
r+ItPP1zS1Pi87Ki+xZ6FEfmdRlDbBoaVn79OhnzZwr+YNwRd+SE6c5NZ68UPVJQIeybsx96hJNj
gtQ9oDdenkrLuDR3DvIvkHSgwf4Q6jGDDvX5GDRVYRFce3ygG7t/piuBe3vOfj+7Nf7cPZWVVzd1
Dbus0D3w8339e286Dyi4I0jDllHEwOuEH2bNNTwj+9Z8XXervvclJRerDFg59DuiiVpfT8VkGVjm
Kvv1kjNGcek45WDxoylXDH8WA5jh2O0dLIs0CtWz2hk3PRXHTK1R8DxGWIjFcZwJC7k/pPvUeU5T
CJLakLoHwlB5pQpzmSUi7QiP9nLDDTUQTyxPxFNZX6LGxdHsq2FpyHOGHY/MckoQeRQj2n04DtLv
OaN6hBLVJ8dSUkW4NSqIPJjtLpbLekSsuaETGzmBCuVh9sIKOTywNYVuZ8cL/XB0QgDzHApJshYW
GcK694dBQrQfgEJt0CPyqyDAHfm0YJk4lS2qMhDvFhsW+wT4sUUokkYnnSwI4xi0h7uNjW0aVi74
YfSZ8qo38+NKw4qUgwz9jGJgIaxE3qt8+9WxIuEsSjvHO61dYpJoXEUpZjPR9AS6o6i6EFSZazko
Gqov5d1ovt2PeLwxmO9Q1e6DL31tmTvNSYkn4K5qW51YdMnoryWiCCfSqhC+7+RpXWiJn6F5Mr8c
FDu819Qu4a3D6SmfY01k65pZj/MOOHEt9IzPiOtwl77rMJtP/KqwwxDdFSD4DP28809N5EzhMRGC
LSMKd86A9rw0WveRIaH+wZ6WzMuERUQPAss36yeoVSPcAscG0RtDorqjj1Wen1FNKF2sEresJ2ER
Y2YLWWCUuCxroRSmdT6sPWMV9ILxDqWyGL0O2MWWRjne0bqqMH858Gea4kh8I2MbllNGmquL5GgA
/+ed/ohIxHIXJxHhGea+5WzWbxFRib2iNlJGT0wuVzsttDeLIRigluu86sa2PwQ2bEOmg03RdHKo
bWDK/P/zvWSp+6mRBAzXO5bvtE9PlGYpV7qijux2tXuNLVWujbni8ihvX7YIoHqATQwET5MVju8f
1Mi7nohNNp9OhG5gSTFlrTXeekNtrm+v26kX0PJ5+YXO+0j1zHaEssvH7zRL5Pm35xShK5sv5tHW
oPjpfwjJosW34alZstWmUYUxIq3EHacI1zuTbN6hl9ux8ZemskGsV5xWsx8znE8r9ppuuqmFgqDQ
n7WIWb5dS/ffQp5l5+koZidc4YPI/x4otzVpHTMdGtUrezFkxEQXlzIShHOgAGWlJ2AG3cWAjpuX
yQxsjqiWfduiT2kmBP9JcZfyfojC6WtREdstCDwTeq4uNm8xWeR1s5Xmn4WBSVHl95h17DWHy6Ls
YhUSu76rGZ/StsPic+bWesYoYhmPFmfh21vAH1epKFZYX+CkhkqUBeXRlDfi3UTiUqv0CwCMuStE
4LHgpq3p+2Cx57Szn3LG7X7/yowW37ltfWMWOH7qh+vhDCbDuxlW6CzoSN/EsnttSWjQIIOw/QCD
csq+ArrueTyG65UdNYH2HMOraBAH2hzW5fGZWooE4A2/O7CF0t1f/0ep7kx2VvivE7mJxhYYHO7c
F9Gtw+SM2uvod8x8Rlf2OIMAunwsHi9s7urHNdiHxMnmJPpBymBYgm9H9G3CogjCsH9mujuzdHz6
d2ML2l7hwTMRHRnLIR2pKiuUwLy+/Brc3lNyuVbo0iy8WaFGV4wumEPpzufmRK6RQcMhN4KONCgJ
cT1qOEsypHDoZnPPmu/l4O+wWcyUcp6cwP21KowR7H39+jn8oUlFUJg98+h6XnP6GQ1AijKGRBc2
2xmC7imUqaQg/ln4u8oSExgxPEdIUp7h5rYiLvwk/UHx1p26/PLMYbw3n4RY9YleD/UsDQ8AuTD1
5dLud4eK7z0I3La114WNK1d+uMza5MRTcrCjfj7RQ8G2cADvVUPJvUqP9g5EmgScONXe1w5jyueF
lyKmmD5B5QMZxbWZ00n+m72Q+i13Bs01jqj1C3xOwPMXD+J0+fb/IP1yZLpI511b4b51F/GWI+nL
8POYg+1rL7T9ATJs1bhfzUmYsNFar9hKCiTvZSNTJHP9uWPSL9UHMVLTJxRSnTVqKWsrref4qJFJ
XbKZs2MORw8yCuaiygBX+57T6TKXko7YXVOI01LgArZn4L3xEIIDOMo0KrtJI8BSa3ygeBqXVGos
KZMTWfLJh2tTPw6jqp1HAnAKxNhY4n5JlFvwJPJEeTRgjXO8QhqjXrFvgviDKW+Xprd4xt0VYyKY
5mFygAQwr2PicTeT9d1l7KezMjB1tMQEbJJTKkJyF5kbYoCHoUbWl9eEwQum4KPtVWa76jRjSDO7
KKs+5oJSmzc3OMB0poUJU/E49rFFy8bwgjyRZBVVsqQHuAvcRxMtDRaR1W+9rdwlNzBNQe7FzOd5
eieBrGtlI573MVds+UuYjr4DdqY3DdANyoAbbeGfXxV5LOkJLol4f8jneNew3amwnx4IqrnHb2Th
vAlUoxi7ApIEk7J889ILkdjaios5M7UxOGDxvU8jfbX52J1S7i0K6+mT2jqdFWl6j7uT9xQ0eFUa
SLjqfubyldPlSVfKksk935xP27AfHesOdSPkTdKMJkzeCVj19IDj2tPCwh6kj/9Vm6ZjTbJno/wU
+w6cQ+qlfR5IL/UdX00FVqQrlY5u8kOtY+MwTYaEcOgZ6r/sD61rjAAVUvpUqSKwKUyhFmetzHqu
dmopl4pu3NTs8a8hZKfMXUHEO8J/wSxV35PKxKIYhndZ79GOgHYMyjMWhYYiZQrrH3qQe1jxYH7J
oows1OmArr8nZ86FwBIwQZWTjHnsh22aNjKQLm4eedDZZmkGlvy9K8eYY9cZS0R6Gusiiax5Pd3b
PMcOTpRtVCvwyp4tmx3mTGF7pRHbCSoAZKyDfuw+IksqPq0G3PiIMKBlOPrCNpT1rGEEYSS1lMkM
GMmKA5TcJXvJVQYC1uCGg/iw0ohu8gxD7x6FAcead/lBY4TKvKj1z176juz6r7ZacBz317dfDuMi
s/0zJWu/4PO4ptVCmApPYFEdsmqBnXw3lttxY225p608zj79OzkHYq7RarbGFyxiRPVyInVyw5pE
xmhMEnyJ1quJECQtTStSAxKUBKs0NWE67aMOLhiVihPbM9oPD122Wr0e52kP1r4jW4u7YWyu/MO5
youNnXRq5FgyyNSgCFzMR5y+sCDTKP3THDzesSHsNoIMhnfpBOvMwxwfYBTCyJcp86if8yIiO6ki
vwsnzB3D+XmOOCintKpiHxzd+X1fEuQikgDkfZCMv2ijBZwFRJO8t0R2f3EBFNxjoN9ibgqFLfd+
spIseq1oAdkmd8yotB2Vxtd0mhuUM+6CGQkkrExCNeBObh2j9jtu/niIVPcilIa6M6/Jgb0K3xg0
+cke2iq6IYxqvMZo5ex4JeWpi1nwSX5CxIMHcx00UX094e+WfmY/J+Hq9aAJid2zPf6xrn1CvFeP
eQobuzRI2ZSRxiQjbozFU51MysZ+ajEF6RFsrttHFNw2H69/E7VDLpm5ZmJzyY/TXFS+6+mni3sE
rSpxU4FBCyNtyv0XOyEAZkaCG6QNGN2pnO4dKoOa4DWxg+MiRxL8uv8xe2mWzVj/cbFfaoxO5d43
XC1q6mOQAdRX13sL5JQ7g72LKNkdO4425yd46czUqVYOB71wtbljhcjOs6Kd1z6dDTSSdCys53a6
sDL90LxMCY1sY2Sd1v86vjbxMPnDGGaOxHTVKH95BWo3OFGiKp7ymfwCwCNpFpfE+5oRpDt33ABZ
tuc4oq0VhSsc0L3HRatHsL8V1N0ToLWL4ODLRXSSl89JdwmqZND9k6EF7Os85Gh/iI64w2Pj8zBS
ceITHIUiWzKmHTeDcua5Xm/tDowDE4u4Hi86VawpFP2aqwLnFQrTAYncfTqC0A+DZikrHNLgULI+
xKSAXTHgQBCM6iKu/ziFNtz4G/pouG2zC/2dGwlHdGAjJyFMjrLZKoYSDcf9BLWA5QFTSlzW4eQ0
vFKKXYc1J2DhYIwHgYvqzo0qvBQcHRY8JGV+ZBkXMPpO2jAda7jwvoH3KPKY8qfcKDZ2/33l3ftS
bB/FG8LNuRhyVJuKARN5srklI3kiKM1nCyFgkf+uVyifNayIHcz6ojmfUwQaCv0PYr2MipyUbDa3
vhkSGzn2YSY4lxLyP9+p72QqhFya8qRfaIuYeRtRHEhXyU9TyEEf2X4tDcV/i0YTr7NHkQM22FKR
7zffWvpl/DAgqMlahvagzNybU5Usu38HSXsCPZ0RH4MkzxHtlNRehIYzoORgEr0ZWwE7xQCooVf0
HU/CldR0G7eHhdjrzeW/Ge73W/fVqXVlQcqB5lDiXyTnONambrV1HPewIjnQCwn8vQeIkpgOlz8T
jzdJxly/uCyFBXE8XksPcKJwCSwYi43wrGi3bTsaIDveDH2KBVRSGYi/5bt62UzuDH7xEI7x6jCK
fsMprJubbbt36+795nRvroZ4U6xf1BKtguhpS+iBG5yPtYQ9eCgKkLIxSoCk7tyCpW6zRjVBC/DW
shK/6W3kqK23E2kMbq1oFndfz2yyF9Lg7AkVbhLZx2wEY89S5nDhhdti4D9oeS8vluJE8PcWnC+c
Rc47b4MigXfqNpgiS61IkEc/4BKdxZV18yQmdwohhQfEKWZcNVqpwB6+ohvBTRf7t0cZnuZypcdB
VFba8nDjAzu7EOAAn1p1acyaXD/VrB56Eg1R53jfDbgpc964qS8oErOkwUyr8lfR4sQMpkL8KW4Y
cfV+bzS+4pRCwlmAvKrzPoqPGsGXogCMbUXglhZ6nOf+L4QO/Ugk52lzOrH8W7RR98pRhm+GTYXv
zA8I3sJPxsXNbHqSlhPseSHc9cUyY/pPEYVHWGr7cPGvV8v8WV0+mMtaNW/P6UECybmna6HpiT+q
OUmlV8aE77OXD6UvAF5HRb06k3Z+boi3rkrK76cIRdImK11uGdZBj6hx4y5L9DN8mVoukjA/o6lh
naPWOrpAm+JfsJFu+n1OS6wsdn3Hn3iJDvgsnlntZwne06A79J6HLlVTi91PMv+wBoHkYUyjpFbb
x7x3WWVCBl92IKVR33cAzguuClICvGMlKNQKOjxm6QWajNCLwhW5ncNG7ll9HpNnZNWP6CIRMu7R
T8T8rJormKHZUKGQNFF60aMbKU+pqLbq/pFk3IED/UGhVWhp87XNC+iG+tkK2pKdW9GuNQtQ6Qsa
FjOk4ssFgzta2mTmI+kxdiw/51ea3nZdbiAxI+DMBjKw/hmrk+FVqgyuABSuSfZUdMLjk3gvKcnA
hUtqZutphX7IMzeJyq8OykxaLBRyw/aU9Dy187W5ZAQazOuNvEjORcilugNHzlDPqD/Ec2pdhcYm
Csumcxf9K0DP1zVjMxQaOUTkpMPbXUvZzPONv1XvMJ3HgHLOy5J7WEUz39tZMuXlxqJoWQm/48dc
uFqUIQa3GI+NsLaQNRkbp6W8v8OWfdXVm8e0pN3v9NtQIHJXNl+fckBDAlezEy/RxGeY8rNcdKzF
6ZERfjxzG5aVXxrh4s5ph+RXBf0vj1EaEszbjg46BosaFndzw/4lPfzJti6Pxho83jDYYlowvI2H
HGIfVkPLJOB+wf46fa5U+VQOFqj2RtA3BujVzH87r0uORQnOwjvBydjAcZqI5PuMbuNy8szQ0Zcz
yfaKWqKJtUJIWw1IEUAPukyVrx++D/H95OLwIyU0E0dhoookMP1cW4XXGrNiUjWw306T1+quVLmi
+Sd+pQ+DAMT/srrKpVgApBFaMXnMLAwyUlHygSagydbHXQ6Bj8KT0QLDxtCFd/wXEp9vj2962H7J
Uvuy3xE6xQlJnRwT5tQiJcpbCX+hSZBt4JGXgnXgkvEEyt36px6zDZUTznTSDsFtnt6feDXe8YXy
9Zi1l9g6zx5OnCSoIJsHWvLooir8t+6/XpWKGCTizDjVU3nJHQy3lVbmHbjbejozDgf/m5SQ+yN8
ELkt1egoJWbe+fiZqRIKDzxor5aVO3G9HlN498ZuxcvsTZScczhSTJ25CbcVpZy6CesFyHsI+ybC
xVBVPnvCtrEmO+F/cs29pSXxY7sveV8TFx+y0CM1Mi0LatjPxh4/K7VRGAZ4eJVakxOQpLvEE3fz
uqjqZxcu3HhxXYpDseJ9qmP1tU/BevnnPru9Nt7VVtcEq+RIlXYG0J3EhRwXMr+OjuY5DIi7FPw5
oVR8opPZ4ZobNBsY+pw5v574i3uXrlHxzLKiKdv36yRmAkHxkFppDW8djKXVF2lwBGt5YJ4m2vKC
XqlisZtDFAGRQTFJkY4Wrg3zCXx5Gg4bc/Ff2mc6LDQ6ihHlVmyZHUDKKbD7BWrMMQBQ57CCES+w
f/RAh5iPQvfLbuhL+T/C8i02WuRpE89COJty+rXZU8YhKkKZRaojb7HGUQto/vT7fMR3ohXJDKKM
DQrDrK6NFA7PlrjKEnSWRvyYcK4Zi3UeYs5HZtF4gMfjzI2NVV0zGfVkG4/LUaYT/L8XeM6oyI4g
bfrQwBSHG1IUsvr2oKbkZg9IZAifNKpWc1NF95imwQNXkmh+ZrzNg7/Y1uQVm7HmZyAT4RXflu8V
Ljo2qFJSRKhojivQt6pFacTezofQK9Jc1Yba8LatSY/dJ86+8slKpPasUe2e1YaOReZRxcIH7xTK
QKUuTQjRACPB5IMWF8/qXnW1pH7Y/yD6t8E2DHZKTCAzYpxkmWEmKo5/qXeyZsmLKZGUW05hmnBo
HcwJNfCLB6ljj31XUAZQicRQkY9xgpC+QXx0EhMbU2nBhCyjhZ7+Tj20eA5fJn4YHzQ7v07cQpLX
hRuztEfo8v2l48BxUD75aetsYNJQsP5SdIbewwyqVUaCdFrl9YhI7jY2szUqVvTfKsYdrbRArvef
At990/Qnwa8qs/RqWeDD1p2pfYmGw6YLBamKrRpB3RCQ/CC9ycvSxgf/RjDeGH2LhxVACQ8EBcaA
OdCPyAqIMhg73dspoLPeQ+nlSevfNDHMSHyz8YSKnwcfLlc8TfHrvCCAsugDjqOT1dYfaBRuX6/G
rkvHPyjAVtDuunf5Zw1cVR1D+P/fgqbXDW00xTmMi2lP+9tDW0dFPnYyNNReIceuJKdGF77SGfSp
CLDfReU/BDRIOM3S4O9vHQnngJ6cdSWVkWUIwzyiLXMofJOBvavgee7JyPSBXilxFvWU6KOh5AsV
HlPY8ntSmjcktGHdDTXVB5uZ4p+EyuPMntJkYxnd/VOMPSOvCd+/7IhVMwKsVWLzWtgmv2vdlfLz
MENE8aIBXljoBkr2HwCMjif06E9Mn2hrOPHQOOUmr4BV5ODl58V2VrHiLf7ZpsuCjl1yFNLp99bj
Ghycuq1qUujgCwfxezmtLQHyfFvBPiefcDBbacIo8RJ+3rbbnMa572IHvgtmLQqr8SJnK3H3XrUS
FUOKeBA6AsHlZ+PbtRWFPJQlJlmOXlXITtYJLpWnYb0otrSPzJwkkKl8fmMZ7HLDghC41viiOuqm
Y56J3dgIYpuG7gZGqC0QPJoy7NM3C8NDTCXJwDDfWKAcga9/hvhfT7SX5xas8R963dl0+3T/uW2p
N/BzffjdUnIU5RFBJmBAWK+ZOBDdwPSg8uxVyj08pNrEDmCqXi5pEXeVWV/38CJmqriHX5pc0dyu
Lt3na+T+ln0MxuTxV8tx+MaHHNDNZ25ZRcARwO5rbtnBczyqDBN7uJ6ywnutOzgvLzpb8kpmTJJW
xd/8YQJjHU6jNoFeaOcicN1HujEZIo2RG+pWclSullbMAQxfSGmb5FZV4GgSuwhWkQRWona6eC2s
3CBW+vGH2MFCHIZGAthUJuOm82p2/nTSgE+eJZJUfkQbgcKPeXotn72Quo4tlF3dx51Yg3SVcmAC
IDO9vMhLOkzo9VvX2cgnPXAfNCCy2JaH3bx1ZZobqe24pPzYbVpRdAVzILEYJ4ZMk9e4OZFAUnSz
4KZCFNk3kqtJBJdAo+JrJtHltsJ4L+qgC9eXWDcLt7Gucmt68EZCIb5fjLiYnXjIeS6uLo6+P5b5
nGgI+HO9EkrvT5u2suUguw6RWaFFYwFrJsETNS5VQs8SfbBPM+a5I2ZjiiDPNVAGMxF5KpZAOY2n
MJg11KiooDEaKdI0in/2RxmzLQcgc7zQvi7qFO9UBjheY0mmbHsTOAca0/OUGTIPlxonQUPq7Jly
CqGqhQHCtI6GPph/GEPtUjEY0xUWJBfGzPjTGYH1Aabm4Lsg3/SNgBbZnzPwlDZSlwZQTEL4bV3k
Ieu/xIE/VUs7J8JrefI0FSASWWvvW9O5LHZft4Xa49+4UQMS7xqpFy9B84Hs6oHsZX8/nnNnOvHd
9rYVacD4eCNUYEqP4UP+PifPXkiDJD7fewe6qWZQim63pVsWi5QcJ858xzgkdMRxbBGql2wiAlk6
yRI+dGdEc64ZfNjqkx571ys93HlzQ+QX7smsXGj/AQvn8AMEUfcIAlRQvPNeESHg3/kBmRjQXCOd
auSHszuXrSiO7QhX2cNOfrCIpj5msdM/Cn41yJzQWF9UodP8lNWcqDVBQyjahjRxIxpfhn3BzVkO
u2RNlszEIzZr0rxruAw7fywT8crJRTaGsaEaMnG6wWNvCbbAYqtbi8lP7MzOeNhTx/ued3lcHpnV
BZa8bAiHjeq9i9/dVlRDRTGq3NBqyE1vTodlV62ktGJFCo72mAe3twh4Sfcq59Iz/1vzbLDXeiJ5
0VLV+TXsNw06aa6+Y+a8nwjauuj2yJS1fnrR0BHnjdSqDAJ3yHioJ1I4u4rVBWSiOt27AORL1D9k
lIVzP1rbkX7drbViwa16bSdN5vmO0jpUqgVbfEjlxuobesaW7lVMV6zAvkCHktFxM3C9Z8dBZ3e5
lbqcVL1qgDsaweML6YDhuNJ+3SyJCGVeXWg+qUYfmS4NUipVhUZVh0Lk5EdhKh915DKuG4httfgQ
s5kOYkHnjFS2mkDFNRpHqKdyvdI0BN3T7Fqz6+TNKoQHw+lHLB32B7kxAgBqmDXOgRTD4gl8j+BK
3BJaAt3ArBcqAUBFa3v0Qsha5l6trKhCHgU8kPTrwBlPLOTn1b/GVog5BkSYpUY+FW4o/7EWHDN7
P15VBf+kx0sZOqpEiOzjRe0325G50PhAZbsSwBd2VySSzJRthppuruEOizjgTm4KS/O59KFbm9F2
KRmxQWhVaikBVcUTV6CF2SSXJggsP+pAdsfXP3SIZ0sdNtieEhVsHg/g62Ct3ObKeo4p0Upy1jcb
DWx95mtDS7j0WZRHq2gEa2DSCZi7ogqltlf88IivsXjdAu4EdzpIc5lDK4Rt8LoDtqgayDaJvQs+
J4Xz5U07bvaoUlsXltweI2lBX3TCYHAI1hvxUIhPbB0mORPQP9nPBTuR5hBvK2yL0fHRaPt3F9G4
Uf9AvL2Z0VUUGOgL/lL/zf8MEQMlLOoNYMPZ7PCZ73RxShbM32TH2xZkFnEDi/6vlzjRG+cpb+Z7
9ePm8OSOOhWZb0wJUaleRaUms/9t4NrN3R/04aNGmdejTMR+uYZNltzhqC6ptorzdqbOtRHBOFNl
ibyTJ6Wg4ieRtpyHgHCOkksVF0kOufebYxubFttu6kF+BXFKYs0+97cfDSaUImCjjjJp5FUZfyho
7CAlCHz1eacfwvDuDXyT+jZGTmpg1lpbcY594P6nWdDSMQHEBiGiTtFnZA9nEquFNIWi2SbZTBv6
NvyfdnHojJ8f1J79TFssaZ0SyDcLgIBMZVNkzlggH7d8QtcYtEVosJcClX612OGxrzwGeQxmX39X
9sv1pV0W5beq8LbtLeVJNn2MbnPW6Wh8atnTKPHllhQGmFOFOWYf+Z4+p3XWE3q4Ym3VnMlAehiD
VZzfZyJTxDT1QVjl6LMU50DdvNjAM30u5A97iWiJWYDQDagCZHWn3sP8HcE5Jng4CjhgEikDb75s
cetlD3Bw/QGtyHkNsl5VeTUdt+ZeHVueQbOO+EFZEojD5V2vAZLi96V0PaXzqmdyqwXjeWDYqT3f
1LoSBJE/hgHwesRggOGmmUduv8Gd+caNkNTRv84Zhm9QnexROqdAM9k+0zOuHg3xJyQh9N1mYJj4
2SRA4WD7u4T7M313C7WSDYd5jovH4nazgst5mFWDaGsX8wVZfw4CczpkNARCpD3ZcAxiyLcGzXbb
yF7EyUX7x3jghrkiq++A3Dhlrnw58cmrYYIbWKxWNAXyzNdEvMrrQgEeAv9j8MKWn1VlICxxdlaf
Yvvlb7QHx/OxGOa4jA22dF+0AsWHmMPi7z8U/TAphfPhVg4W5woEV6c4V3KZR3/FZZVFIzqL4Pxd
M9kHbLHfn6MIUlwV8FQlW2KqFlu8HY9NKBefphsJd0wfnJYfWHSFZzofEOne11DqWmCFAA+1XNUz
bjpinueGNIQPXlZpqYQZpvLvePEumRaNrSK88/KqJb/Pkv1VB19dtsVTDkjlD/xDPlnTLP1eENyZ
jy1WKd+lc+IFTDlflJzucdiNOWbj80IO8fqLhHwPsmEzC30STzajtTGU/3diN47aBAcLGC9xEI2X
znh80cZUAo1P14SRYS8GEIJuKX0athUUJph5fTOLtXCNTlbOZkT4CfPhzcfiEnDsobD3S+B4pTRO
hQp9cfFlUy+ClqZrpJWRiYom76tClaGyraZ1fpjJ/YHbOjUA0/N5vSAcQbIRrsgbnRQAmckpKF70
mu1Bp3IAoDRhwtrKimSBITLVdnYEmeKBs4pMA2o1nUFESiM+qc9/ueM/Mrn6XzuHelCA5adN4/NB
xITpPpV4Tg9CS1PtGinrWEr2A492nms36Hfa5zMtgCUTF0U6bPFMc5KEdKm+pYsqolj6Wss9GjPQ
sZN7Lrjv7or2l5vPOueQKaOcLq7v3M4Xteux2nGBJmXNRtgxvy/ClINrzWR2QAIe4DRT2N9JLoRV
jb5T30qvxGo/23KtwdpGP9kWPcImwyH9q4Ke6l537x9Un/q/4RatJ9508eoVFgS34b6TPoYrPcny
GXJDWgLJHacxaGQsiQ6v9/UvSdpUv0QRMIDcYN5d8vv3eaIFbSe1kzmuDuVopkD77jzD5VPvA39A
wbKhWGMziH7LvmgJo+j15x7VnzobSFMkcm/yVThvmHMy6cf7htBWaULaDOuT7XjoCxsiRo5oO5dB
cEHyLNR4o+2V/bjJk+58wiswMZ6oxAl2p3looNwe6UDl6zOAJwFC0ork5aUIUjtF7IfJUawq9UCN
zwtpdK6TXQAYBpugz44BKr5qQ7cBIx6QER+MpjaARc7ka1s4NMUi7iUwifvH0EGA6CwA3Z4qzRdi
RXBCVOLpv6m3ZH8G/xbPsCjKcuE8hTGkLLwa+I/oxQZMO0psto74oIvFJ0ll7FXEI1ItrFT5d3WC
CEbA53DdqysQ5dtoji2tSasCXfLjgOA6+q+HgLWAjs9j3tR/aSs38bN3MsBGYrRkyCijRO998Zz9
qRRlkHuqmfmXbnUhhYFXpTC71zBcW/SgLSdUQY1p5D17KQzRxKZpD+aKFjIiYCKWTrOHrt1sGD6L
VGfbmzNabcPRt6oe8IsSvOBSonPdFgXEy/N6nHSIjqu3qHjblh773YtV1l7Jos6HgNj3wctpzITV
wKuFxRKiflHJbcZ/q0xolzYKUy/jgvnMlfnG7WZLJbzC9hXkKFMcISBwNXrLfxuUYMrp2amwFCHn
6hFRtvTb3aBVP/iVOjYQQ6GdgtgLDtgy1wvkpmseFtVOSf9Vo4P57WMjMtmfPduqrGu5DgBOpMOT
egaX/GwTspightVe/UvGbg8i/K8znEIUxez1kuC4tgOM9fy/aHJyIkg6zNuqbc+1VtIb+Bpo02jz
ok0ZaezBDyjnhUV/K3WaI3E04fDWXK64hMXvYt+tSpI8Sd/q2UUz7s8Nlshxjew4CT0LAW0Qhbfx
DWFv+42DVzMcBadNhvLXyUKOBmgl02TMnnJpZJY85U7I/gpOM2Zh6hzdgew7y+A7nkaDvVz3w/Xg
OOKXas5IXZO+zjoKi0DwkmV8EPrS++/HVws4zU3rG6151ChY1Jl94+5VqkYZMNBGFHad393qoffZ
YqqbypDJ0iKkwuXP3U4lKPkR1GMYTwMU7yOFUn/Qb4LxTVyBPfDZPEiaH/UAUlZBcx8SU8Cuh6ep
jCGmdpaDlXuS5SBw8+XPmXdD2zVZ+Drp6Aj5sMUekb+qelNc9AAofyJ+jIITEEHzvY05m0ggAEQv
BpYHamhcHYNcVXGOrZdwp/7iNYj/OUT5QVkBgA1TOgUBbE1VZOI2gBpkXGIC5bkSFle4nxB7Dx2g
g3ry+nvPena7nw+f4qmV6UcN1oJ63Ah8W6k3DZOV6vogCrGj7IO1tp2avmoTqEyJtJwS5O4vYEkO
h47LVeWVHTqGXIGv3/ByOjFCNmzOhztI7EPNleA7y6pr/UBo2Ruw8aOCYnBAkvDQtLseqIm8+76q
1z+N49d6TqpbXEIwxbzaYjSkpRiQHhYFShi3qwjLPiZ1qCp+5vEd7xVXDRueXoYk1xoOD+VZxHv2
cLCofHparTqWk1RrAm28CXULa3Bkh8n16uS++X+wiIrTsx6HOWIM4hoa1WOAbnmfZD5tHiO46H0r
GaUD6q1gqHA12kH6WARZ654qXpJhOTP2MdSACapQ1zI23hSIy01HMPKoj1I39OGkiccgxUMXKPLO
RqJc5rIg0X9JyRz3sPEZ4c0xQ5tjjkolhw4tdlLDBoPqmj9zsl4x5Riaay+EfDGUlje4yE3YZfBk
EVQBhWSkGjhfwzT3t5Jma/LWpuj+8WKbcgXjUjBNdfAiccZrZ17PpjZwA2GtOWpaNf1bkr1Ka9Te
II4xLlzx02BI6wO8LZEKTZLsRzpHuZbIGQiV9KZXZfrO3+7QJvGuP/WUjzVWCIpFzgeSAx5uKxAK
LDBxjmFzy6ZyVnhc3nsLoGygjINo+JaxwmeKIFkdCMGr4pyjVUuHQ0+qTc/s2YvvBZBQ/Z3n0vpD
yyMwQ0JeVeI9bXuUehR77EMOvYaL9rJYThPFvLGGlWafVSr/1q257P/8WZVIiJCPr4f77SQ6ZS0X
o6c7uBr0zfiLJFhvhHJDbCRo8ju6Jqo6E605sYugF+PgNvDRjAxo89H+AF64X2OxpFVObRXMWr+d
iGK3/CTiNEzQW1vXJZgBYWhPLW8BCHXIsHhDBWe4p5Wn7M6aEU7TtslExSCO9EU+P68G+3QazIYr
hkyC58aRSzIHfZvQ/rQ0/K/DiuPNmu0lZ9kghiPAcgKze3bFLfDVIfccLY+yfrq0AMUYap1RPQ8p
yUy0WJDOOL9uCuB5oqzz5bg8fqdzYH4m5OTEnp/ChC+qlYdkjUCxYTjMxJWFjDVlSC67IkbYAM6W
5OxIjOakCcQTUZYpFyR+L0pnV9EmtxeZfoIlyiNwIvryCOD2kKu+0lEZXX3Qvy0Cepw8R4Q3tKRV
5PI4YzRw1HA6mwmScVVW+BWzr1YeTB0c6+7jJxb+8OLYVh382xluE7HUPw1Kl/kg3kO8Sx26GhT3
nKeIqdzFvIYJGOPx3TIIe8HJE4A50x/it98oWtMJmsiG8xk1SRiDtJ9dgE5y0cZm/cwZH3DepWtk
flWiZt8AbeBgufHms4RSov+6W58HCeh9eid30l5IpYi/G/R1+Vf8jvuDM67YOWeLHRQ4rg5m9jY8
/rqPYnW+P65cnxcTIsIjQ48y3QpZ41LreF0BHu2VdEw9XMi7/Vi6ZZ8HNxWnQMRjY+GM3J84Lhlo
4NlW7S0dReVslfp9f8E/Us6B26wFVdBA3Lj86rHv+XbWnh6UwI3bQNKbxlKCGz7mXCdJfLbNjlOu
G9SkZrbkP105rIA/eVRiYbQpebDEzxSmV/ThUJpI0iSVH2fwChKUx5gpt8WLjWfhx3T2jVlQVvcR
GidaPqA4Okjjf5W90XTrh1zhRhxATdhwPheDb0/fQ7IHjkdPxTw7CLfUortSLquW+mfwzwUM0rZ+
zfB1Ps2I/iSVsfhyf3Ed0xwt7bskiQ/E6PLpEsJOEgal161xM8dXxQdF5+h15EDkRPg6i4ogEwvX
EQXRfVEcOyFMsNxThAiFQkVYZKPTYKDRkpWI6mdWpyq7HwyFCoKWMtCV3qOryk/lfUKyRWT+4XIu
39xdAyXj6XvTOV6AQ+l2JpVAr0cYpM62eBg4TFlGx1HBMsqZK2tkuQFyaQwSAC2f8z3zUudKkPdq
grtwheWTgx7toMkY4czp+UGPoCZqPVyRlttCODqj10MaGgp3H5sJgyFjUcuai4WSChU5efBALgGc
gLe9UMPCk3lArUyaQEGrC5CfcXcGbabih0rp4h4bSKXjfdAhJ5tKpAmszutqbbkOwkVV09d9ueIm
QjbEfwkP6GGTlXoFC78OizqwqzRq3m2trWFmontf94NdWOb16CD2y9H8CxKwMnGeHNhncje4FULX
lKHapiInyfo0OZ39oNPROreYulQgbQkny+vYGEAYKmyUJx2NcHlZGt3ZDQ3oBK95WCOf9vV3XV1s
rPF1f1V43MPNEqMaF2QzyHh4fNe5wrG6mS/0GtcUgfFadpLpfQkHPD4+Z6Q+jNsn5crA/HLesvEV
4eVN9/bwhyhBRr4wkbvBC0eBTxj7ePljikDnmYb3dUj/B2opveiF23FbDIzJCLAdW9CQXzhSIEG5
fJlarw4tZ96H6PjAQgK7VBBjKOaLrKoA2Nq6fnEChVoEOAHwM6i7EMDYFXA/57sgHSnt2WVFiZ20
jxjwzLKBRRceRDRaE29Z5+CzTJUjqDoYtVD+AHLUu0LmNXDY3Pw89uMblmUs9uxcLCmTElXgajBH
RV6Bj5pKefLIO5Z+s2oTgIXVDY1AYN9mKtM1v6CFVeTR8YyQzwMUt58ZJjffjkwGvPL/5mYZqO9F
8qlFcaB+pCiobHvrIMHuMzdaA0DzhQvyqyX0VJDsCMyb0v+lEpuFXkYsxJXXo1iZJUswaQCQSRGQ
aeEaO7pfbbEGISk5isziWaJFlc0ZA8fF06rmpsx/71AS+vHl0IwMwV/Z/8D6Gh1qSHC202cET1Vu
NRN7XXkc+cigCnqzc3m2Dg9Uxh9MILf+VgpBtiBSoAbvQje+nb99YrRBgJ8q9p4Ylv4aUzVFzX8y
N2A3G3o4fz+Sl5mTZPcoLnOKLIJf41Fc6BOQDKpPGcuaaL156ntzzBaTjmW8AUD/nIKqL9BvhFdf
/pXpl6i1+tY06ohDH50TyMENvREQ2gyQIuTt8wBsgEsZdiFIQ2A2mVqs5cx+8Fd/JHA11U1+0jpK
9eIZVmAkUqBZ7NKLZJp3C5wnYsjsyfZXAbabtB8X9tQ/h7LFzZLJs1i8T9LhfOxxVuD5numybdZs
6fl/rVzlXa4Ua/5+EvPhvdcg5oFyWEGM6DK9HObV9EtnAw8rVSMhORq5VZehtVE6foqTHA8O72fj
G0VWG+25Tcdvm7GTxXarOwlBlVdM5bq6/IdPc/YsGyiQ2E6Q0h4xBqwmO8o8yiFxq1Rc0HLTMB1e
AEco434F3MgytlkhGrjl4VBdU14fDI9HHbwbQl7rq3bJvWIAITkhvH8sDcOkLWH5E+dx97PxRN6F
EkOrtLuMc4Nz6NbXKNtxppyZNKkas46cfoYuJQZX5P5BWsTENq4H0Xy+/7AvW3KLzIW4eDwHsAMo
9PvPx6QD3nKPeHgiPd13/XbhWXk/O6S48gYSGwfDHVVRcJGgY570ZoMpL3JZ+JWflfc01A+y1Lnt
jbgc7ca5Jvg0P3t3OdZhyAEjjo0VgfK7Oft2wsSff/1lFfYXaTj+VYlkQrb89ILg+6dIuGgB4QNz
/Xyvl60MOpb0sBda4d0bpPzJ7LwmLMCCgof1xjLL/wrnywzE0zUEtyV5eIQXhonxXsmfpWhsKqSP
wZ3b8lSUTkjL5xbSZ0f1arzO13aonmOMQgYhPiUTVC3YIlJ4r5jYj3vC9OmHMhD4qVDlND4TXNX9
8/E2iWQgCFRk48QhJQorsTVJqsZPjhCBI5dUULxpHB1bNewrkG1ZLFMEyd9zhwo4PG4V9OYeiDJi
WNxGAwlDxWT/Wxwg0M9kWQ0qzVBPW+h3PR/d3qY8yjUpQhuSGyMYS5LY9A0E2RxTNVJzrp2Zk4SN
qFcRiIGzEy9VYK8/6ngTSwgEDoWmpntXL7N8/iYEgoNSwThDbFAj5gIVx3zNMuBZeFfC29/79asn
uT91erXLh1XVRCpXeVTidMIQfnSWhivNWXucaGFVzOdcVWLFYLlvkC6aXho22l5NmBWFogPks/JO
saZLISTnVkpTvxFhCwrJ9V9ny9f5urwhjIAOZY/ODbf5ijAZGkanDpiOMD6N8nYjzCWNi5MnO+Pl
5+zXNyV7WNYj81N9UA8xVM+qIUZ5xwokI9mG9w9t3NUT9RofHTwsUbQtdw7hL+p4kXVyovCqh/F8
risoTd3n49RwuQurIYNZkr/4P6ZNVwscTMnHlhpJzjz2TJQPz9L4WxaSzE2mNYSxTdx63+mdGO9l
sa/tJxSWwttg/GQQS1YYCx7U748YFA7me+iUuUC2uXpMhQw/icgJgNfCpklGwTWyCZ0WJiYxCI6i
KBKrp5Y2eJLvZotwmDRLy9LR7xOjaXleyJHIeHXZiVSu6ZN21Vq0N/Ydys8DoK/6+zcqaMLyR2ac
sMrRms7jr67yMj93oYeQQ1SPjFrfAT7cYlnLbweOa9LWAVFxOrXdX03jpZLL46sHUknAbZuKExZW
VntAh7Qj/i4edJWQEIaH/1ODs7NqsJAmoXq7apxQZVzHvaBgoYxgu/13V7FbJpJbWfkilvoEpGxV
feH0y2Ikvld2CkQsYMbK7ZMEK6Fde21OsaelQZ23/GHYp1wVZ6S8pf8kHO1V5zYVphgQvF4fDYac
CGIplFcbVZY+DqgQt2Fw+ZcLuvce1wat7MbxCQAJLWDJ3ejS6+Z7un7nVJlhj9xzRWSU2uwdAYQ5
KkZQAY6s8ok9j8VOplzdenc6a1SB//sB6WR3I+Xh+q41onZSA0w1MflNmC53CNClScPHejjWcGGH
+4FnG4Y+LFMVyR/9W0FepFq2H0djEUPvsS4o+ajOL1KDbn4MZJAKDIrlZLULByDdZe288qApIMzs
SevKCuPfqqOUh3yrjP8juOoS5UWIiTXCZFyYAV4b9BQTi/J8gycHZ1urgOsvgSMkt/eQItM3hNsq
hSPCAukffMtCFgIWkR9gicxTVt87iIMIsFXa8up55lknMcizOUkgt/50N36WTDGFsvoMvaH/AtlG
cscwY26LH4TiLBFX7Hgl+ryUZ1casB6Y1o7FIKx7Ve34KsolsYmARAr5LCyWSu9CG0nUINQClPNS
Mg1YO+vJWbQeA+7xK5nnJQWASs6DFD90MBPoCCwrK2At4xpFhct3kU9on8WUKg4bO+JVSwYSyIg2
WCwRUxJG5j4v+mVIF8n8eDVywEFlnjnqMSINqAlgdwavewxkSfqhaP6GkulvhHVrXgGlxNF1ByKs
gpKvhUPcIPeSvjrSWx9Gmm5jiwbs21C0pwSvDItUbqvVzHhtLQWZ61x65T4hntSErD09Vz7G/2qc
gKG0DLClBTUilqnfMtbGQK3tsTEPu4Qke+mHF+BJU8mhNbauK3aXX+Gix3qiK72MV3nYQD3mcBCV
KRjfZsGKkppeKbdi6vDKnc3K3uQsTMh+siyJwJbMd8/Ml/W/R6zE5AQlooX2UlQUlXCWS7ur6a91
ubu7+00Dh6mf4dzkA7SAn28YQ7b37tSgMseiuFSx2VY9d8dJ3wRWylrepQcajbICMqROqea1E/yU
pzuc9vW38Zfzr7mZpMjlpI8n8O6iRyR4YjW1UN22B0FPypYS/PSzqnREW40iSV1tbZ+7t+ZR6Ark
2cnfPLoreEALDSTix2EaxdA0GpIrTaAxPClDE7Nz4q56/QtqOpgc3FG+3oJUU6xOfUTRV9frh+CU
4/sYAsDN7/H2TzAeQtdg7WUs5hq/vANxqqpZou+bx7+0u370AuSNCx+k2IUzapMtEwWxkiIz51xF
YlHt3lXsQ+Sl8oeyIxWNvAa9EpZbtE/4ZRB31SJjeD3MzlUvqYAwqj3uVzqFjVyHRvXWef+uDxYh
/nAarazhZwhYsgPgvRV0cMRWqsLbWG8IGpiKKxtncMzwi99v4k0MDnmkjoyG55dqJwIjApEkheea
IfH/jFgNGsMVlwZVD8GLumZpGd8NFCCUC3dme6NvMEgJspmRUHM6wss/NoayAIbaNiLakWo8SENl
64fqJz7kPq4ohjksh082pct3ZlJS/R16XFawQ0n6Hij7krJJvwDvRN3vWO+bO8lyN/369gtF5SP3
zKJVgxgTQCCmRFqKlyRhN/lMd7p+B9cQsBsmYw8vHLVKQi65WKNIygRddIDZvXSbhSdNqybcu/UK
yclhYkM7OlKnljodCF1q0aeHVXPizjfgNI8OD1zEOH9+3Ge+HUbNXQoLvAVFwoRL8bNgzH12S46Z
7KYBnKB04QaKS7gcEMZb6/lLv2nfOQIWef/BnrTYCLXt4tAJDJlz9zaz0LwXqzajpoQPTlTxdOnH
694XG5sDF0htjyHewcuUfMpGySisw8EXOd3VV6t0S5yOh00HlM1gtvZAB1+3Rb+DUxHRIxl/32H7
61cz1jJg9Q+8LN1872v9VrCuMuxI5qacp8uoGDE0PjnYVDUC4JajH6y9GkS893PI9hvLz14qyTH7
AYHn6K5ibVs/6wl8+obaPv1+NLvyTClQTIzSpOp+oAiNcnF7hInLKE/TjPWv5n+DXKcKtBQHhdPX
VA27A+3vZN7oa0YSp8hsvvw3hvS1x58Tay4bnnkFpYrm2tStR982gX+1t7L8I7Bzj7T+t86kunok
GFNj62bA8jf94HvvzqBzjfO8fDFQBiNSqVs48ndIrjhko5L7EfPfod1lEzOYo3sf10GqXDWPpS7Y
WmLkuY9z7fAnAmouF4wNXz5EmrzLaQ3921Ip0kOxUjYx1hsrrxq9NjPd9TtPYkOVQvdxgaL38Adh
TchIJ7r+hfP9olT+sZAbDvyPOY7Lb2fN1yUVZyRc8Ea7cmZ6sHEziKquI6z+1FwR4z87IDbMV3NJ
E5vhOMTmj6QNE7pjJWVXweKa2tC1DTJMOIvYUTyaKLOR4lC9Lob7oL3iVuTZFXa4Zq5nWsIRJ+bt
gkrONXHHNCwW3S173c0PbJIM18hT+JDF/Jq9c7rEtgItYrWjCPrxSz/Rnn8rmbUBtqc5jGqXwbD2
bdPCPeLy1fO3x8Ur5NYCnnl2QghWEsNZgqn5PBhmItKePy1ZijCWhwptjYQEmITLcZ62fLIPS2nS
c5tJlsJQzVFEw7vCi7kT31sBZLZ4yS31kxo7AB4zGxSsPGiL019K2geQfO5751nw7xZGDvNJj+E2
PjqClztXCU52oo+CxfVVhwR49lMEGukuAHJX91xfatcnGqW/SmVC9HWhYtZsgUIf/PqDugkjq0qo
7LVBo2VUCvygiiiZIrpXfu2car+pSd7lQNEPckGnzHlNIkP13MUHR6sD8rxeNHG1IfpzAtcfk00R
XJjyuYT4uL7f04A79ihMsVInq3ZQW1jX2AOTVX0jSD42OAhk8fmcNlFypj7I6OYOkjYU4zwzokx0
hy65vkCzCe0e9Z2Vn9oJ00TR7t9h3IKgklcA/4YXfPdg1Eqxzo5ajxt7u7AMq4HgRCc+K11s5DMJ
LfF+ZCfFoegUF4TLyfuyzeaQ72Hu9TXH3HhIqxtmWE6a/UHyC71lvWOp0H8WMlN6vLk9LoyhJ9Y1
nFZcl7Bw202spTHvQ1YNYeGUQtxausR5AuASIriIiPCWzaJv2lECW3bEprLpLwSSJma94euFfK0A
5kQA6da+NxhTk8bo6J/WicGfFeofqg1OXbHEqU0ggOp21cm8Es+X5UsqJugMo+rpE7DK5M3KnB5D
WJVPKPdE3RIW+Bqc9KljfgpVQDLxYWBOQzo4HtER/B+2lyhUNWopxePq/DTUHDsBsi4w/gADv8B0
vAkn1UYFlqxFeH2qvrhfG1uktAV3op1b3yFDGoHmTpbjLJXMRHWe8ga8K1WbTJL/qYeW/m4xAxP4
TBnvHFKNWdoR4LRidbLKct8qButAeMWiTuGeErOKpEq7Q1p9gpeLfFQNZfjb3q0HVmgTdZznGiON
hG4I3hVYmFY2ysay1YYdI7wERO7oxTI8qP2JIi5WbLSSBdAXRh9cownnA9eeY6d8NoLyfQWGMsWn
qUxcNSdtNYSDezqi2IMfx21Wt5OIIqW1oYdthSFfrOE/nstGcM+vjlME6POBQkcKtBfLJjOA+G6Q
waDYzxTSCbA9wLpGUxqJ7wV47OLUo93bSpwtwQSGcTNrDttAlo5OCUAl7YKNYYWUlGgoU2GvIPz4
SDPBeWfyY0K4DFKt9BVzEI+BP5BUk+vCaGu9XxdSJMOfwhwXhtIYWxwFon7j42sWvJKKqnPcuyQy
JO6Fk+JDBD6YVnT+RE67JWU2+J1vQWc7Co6+1U7BTf6235jW8diXWaQLK8/m6dW8cayvpCOO40gL
TXIg6hAB9JRpeODIRP8Z0WtqN5ELbWQaI3hwLVrcLRAf2RM1Kn5FE5DuZ/20NMfutQwFgFYcOeIF
F11s+pRVDE9lMZxZjkYn7GwZLfefZCw09ENUDV/gcHN0uX0L0oIyPCLTcKHFa/waNIo108hpGe3+
YgXUFLEJ2FqimTmCNrykZElymRwNe3uFVVad+OBG0Dpa/7W5He1NNcOCf/iIlFNOmET1qpuoTAm3
vDFBqyIFoi6SC/SEI3lSveiyHLRmEeYevqsaXiP4rVwJgeKd9ilPSv3imQTJ/Is8wpVabLMM60Y7
+1SJXTzmPiQ9FS7Z4r1n8VwU+PuWR5X9xjQK8FSD+g3CY9W5NVNtJkEzRUK/3esPufgobX0UD052
rT+HQJykKzFnZ0QjSYRCpRSt+1S++lVpvdHmBRfSmlJibnVDdusMaTRrtrQ+yqRpd51F8nXJIq8X
XSLg4hYUP5edbaWU/SbkVMp21L4RxfMRr75ZJajrw4IWCIa7IcEajPfJmLnwUfUXLCF3Ty0zcMVI
9pV/hPN5357NJ9DVI6Bin723ERo/3Qsl879kczEgSLWEgKAJid9f7Lbk8Unl2cKlchUfvVvdlB+p
xkeJkpzQPB25Hsi9V0GcxNNGY/LTcQzG6uzHTCWPuYOrikhDGyI0v+kOKLVOUEufczQ6v6HBbzXK
WXZp4cYztDNVP4rmnBA1ky3UJzNpIJMgGNkrxkZcQrkLZ5lH2rre4O9MAek8LEHGCErlwYdVYRWH
dxBRqd7A8hGNjotndE+1Y049HCYrGJUSrVEH0hMbB5nPjnABTJGCPq6DZLv2HyecDfoldc5+zDp9
0/vN+QRCkP2fKzC1ftqN4MwigVPwiHaPmv/LKgCHJNkCrkqxMm4puODcOQEiy14aoSrZ6yueM+Yb
v+Pp9kClxUW7UjaunTcgux/2x8WwqYPvx1Ajtz0M5ydTl/NwmB2lP3q9i3OaFZHryFI21e7l/GNv
sHn+U4tCI008ExoE+3Z47PD/0PUQDMqeKdBnFdeMbDUFE8JMQpMhTDBzTD6Lw3qzCKWgOileY0Lo
8BUezzSmTVDb6NjFggKlZoPcTM5ePk7KhDiov29pHJKxjXIkuSnnmut5NIj55e0Jq5RMuA1hPVgq
9FsJiyrCNCxlhgP8SPgdhAKpCTvFGJcWOVUIgvSTiZFzjczIlAW6LB667FhSvR2uyOpHVcsLlrme
6WKjEcJ9dJ56MxGPwZ0loHRipyInxDV7+X+tdl5lhLU4tfFOMJoFEMtxJ6hxVYwXr1ZV7+l954fi
pi1R8Y2LdrevEyoiDmnsdZZIrncJjA+dpqW0Ac/hvThKpL1j7dz/ehU27cz/lJTYc7H8fJ+pmsUJ
7Q3YgWFZfX+b1Hb8S/csqR8DAwmsEUqv5SE/0t6TXgcsK15cCMfbxli7AxRfgYXu8+JUHDbX5uBh
2ypMHDAeLn29lqUtXVcFykUzMoPp5YYPrk37Tm/BZ9Lx86drdhE/4BsiIWyZmFaagHJ7wu0j2MGd
dU1FlF7IfEaETvuZShE94uI/QxgNUrjGY4XxiygZT6RcINZQ0MiOHmzuHg7K6vnr1nXSai1DDMQR
TubDeZ9yA8IZtPT2XUyj2h3u3eg3zDB3zfygpUg0mY/GVDhEXyklCQhGAeW+ClLYpkPUluoDws4h
8yZg5FjChA3LgU108Yesoobw8G0EA+dn/MT1Lp310om7jGPuQa1k85hhx7SClmXlna1o2Dx3n5pH
6/aBQdJNi0MfDAjjZjyLjU6ACreWZUtPOsdGIh6yzYPVTJSX7SYWqqohPRTJZb6PT3rPZwTjOvSl
Dq+W1Mb/ey2rh8UgWcqPsk7AUzm8iF0FRSGkpmIJfDjDKtkwBUOKSSnp00wY6l3b48bGH3Rx8OkU
Wq2CV+RB7+IjrlRb3oNIwCaJEVzQ+KobFVKs0oo2ouyF97BFLsTFR7OOHKxaFKJoTj2KFrcE4wAk
YiG+UFRE6pefGqAb0cYsu0j3zOwe2NB8x3Pf97o8yU1PSUHhbg8yLFrliHYWJ1ustcKdYBdMhZUr
MpLTZxse2IVXw2xoc+uqiDAg9zrh9jPkbWWxbw4QydC3pTaHcIGfr+HpdfapcDX6h/MxHVKbLyBH
AgPQ67mwXYEDDjdoxxl/UKj++gGLy8L9Z/4nber/RyuzPtqpDO9gi2bV3vWJ3afgvV6igmyA7X8Z
mUZNKm+WE6G2bVGWM2GEgOjlNY5teA594xI6aaYK945XAwMew8SunfGVogZ3y83qbvkDmPXQFWIC
lyI6PSqONfDz9kW8AAlUCGvxdKS2o4xuwLtAvBRMUZh0+GV139LiV9tjNU8gm9HYuoQiaTOYMvKw
truJ48Y2SudqIiq/fJh1FUBBWvFxfqnA28Fi+Ak/SuDjsQEHq0jb0bZaL5XXCegZYh/3d9U7+4ez
7fM7m4Z+HHbzkCEVY46f5TdkNMWj84bIv24MT0lY9eWe+8hjuZJpFmzNjLfqoQU3UDn0rr+gETm+
XFucKTEm9O7QMhaHs8K8F2OeBGbxreZaXBMW5vDldEWHmqwjktB9KoVD6oj1JSXKKaj874CnqgPh
LeOSMQHqlQQpLyP7UdSFL/z4iwj+RHu+nYDjqFVv2iinYNeFuJFnHBwa8GPfbJImcqcTKJSrbrvy
NqJQZ8OIQAy6PjbycOOZ0jNnqJua5W8lqvI/yvlNfvJZDKNSPFSbbNptzYxyew0EILzxSJ9ZtpYM
ejzWVcmGijZwf71igxbzMehuKWfJr5XYuzJwsckIDys+vdYC1iPKF+pxB5RfH8Mfl+DYv8A9ohVa
Y09Za4LLbVhcQT0L0u4xZOGAjEZOOY4nkecq1AAzZBeRd7XOnTc1K62FHxkdVQ+y5/uf7XSaYSb3
g1RiUKIoQxDEhpHE7nnKYCeZF9O+MGeW3vnXbvu3PGnK7PV1Zj6Myghxk92QBnFVmfQFYVThy2LH
luKYGRDZEZxFOy9eneS/aSx32w+4cVXg2Gv4hNKtawln/oFEAvmn8mIkAFjl9ou8EXV+2l/j9vL7
jgOJy6EIRhpVt5DId2Rch+IOQL2h4YvTbsjZtOG0mkeIi5o+uRaw+ZWIJ8CwCT7UTO5NYJUs/4q/
9kQMACokm8JHewGMFmwpiKxPvUKB8odzLieuZ5RtHCAunfGjx1nkYUo5pnhD4AdUDSbFz6h2nH1o
lb0Uv0yqfSEu1TNDTgqq7/ZvHk1h7Bfh9RAG5oaA8NGByiqT2UtH4V9JMGIsrs5k9swvYn4ZySU+
4C2ySYQwC/vIqqpQKsRYHNdS7WCWJjjo56s00RcquvyYek+vWM6glR5yTMh3M9+A9598De7BQmWZ
TdgzQncYSPwgoNs3FbmZ30mv2EY0lx/9MIvl3gb9xCWxB3cDK5YG2ynaaB008ca5Oj60Nt9IoVxM
827l3UbvMPljpGYR3C3sBIFqpo6Wu3kwmydri4u+gyUIai0zysr1IRI+dkp0fZf+uU4oM4idYwB7
MNjVoYcnt7jls/AYjlo6SK6t7OE4M9IK/8+Uk+a/xGMTLeB9CMd3xrKEDkffYVZ8LeJIqPUhjRmc
zM1hUc0XKs5sVNqP+OgaEs3fudMD/lHV+JI/1J8ShhDDwNMOqRbGY2Xae9wXJukDhF1DyFIclKT3
UWFTm7TqePqiZ7DMJZSa9F0RoeBNMnUC8976Q5pMB1EXoO6gRPccAxaGtSUyaGaJ93kCLHcCQ0aG
f22xYFtSTr0y0aDdaP14MYL9UX1/iCN8iObf7Oyai/dYav+upjb98eDKDL3VmiBkeX2M95a6fKBB
DK/JqRgvQ/oQVqeBaNp/ZiLLJJz72c5DnJC0dAW0qQdcgwJJz+9E2uTwcPVZzUpSN2flXDm4HF66
whJlthTh+uJG40Lg2EUfLBdQ0XhPZcL24zRvilqxtDPGUOpez1kyjG6DBeb/ykZ4BV48ix6fMLFM
vvJTqzPFTaSCC7p6Bc+EpGII4dWZSg05puFpnwiLS99jD25EcO3Gh45vvKaPo738ADrootdqLJV3
4Decp22nZLyfzvlcrZGzdqxQEubbH1CfvV0P5hlxLGVTBfjS87bRwvNCg2JrmiX9zvoKHIJI++mq
MLoZ9d6GHKGBff6v6H0dkc+JjwcWsvIuNKU5bwTFRisUAHi4tAJNJDXREfbU+JJRauJ9QPm14RB2
vd/221JaEhWRk1hDmrmMRsYc0lINAGYmZbAcAY2q/RNb42S4gk3L6K0FdGi1FKRfQbydSXWiaQpb
Gphi0nRvEFgy7Tn2yOdym9RoiVjvfh/gYE2UeWWbdCnamdkBGHJ4Ak0/nGxloG5ZMMXXJOWlLvhe
AjUSuf/2fEOduKFKaioyw4LIigfvC/LkQZvVFJIS1xjWYUAEM/IkNkPzbW+Y6CM2vio2KHrUJ1AU
Vc2AUoEbKCIBq4wMr0fbZ5ohVpPX/UXHQu1OUeu+5gVK3nvZkegYmVg1IqRxGJtqKkX7KuFM9x2i
8QhLdmOtcanUqCqksoE0I2uCrtrBkZXKj8Siwh0I2shtADu+gQBtAh7obIf+0BAfJ1S4CVv17/oP
zXNQBlLzpZwzC1yLbElnsS06XX6xjbugjAYGASfnzntLPRIQ46w+oT8e0s0ArCjD+zPAPORENWCs
lEcEVlOIUgDoqufLQorZM7/EP0qI5wlknxUpCSB94pjbykRmL6Wz+1abaR9ab4KSEAJ/FDVYp3SP
wMhyP082oENRm/FO0+vrOZN0BDsgemKOUo7/HSSkvcnOJQQ6b9Em6yR74AIcUaAGfkKY1WzUsGmQ
BEkkIO7xmja9yxQST2mSJIqY+D3PsEOrWsGn+gNS6KDd7hKZ0VP231hC4Htru4dmDPdTtUbY98kp
NA86LsTOJkD+Ae00JXaKPTCzurrqXGzG0UEr5LL+FIkmWdzGHWJ2exxa2oDar2eERJVavjixyk55
RBqROe8Rri8xQMt7BETI/MnJwbI72ganDF6iGOJnhyfPr9nLIjKW/04xRSOkO6Kida4H1DYqK4qq
jsskdEyCBMTsV/HuiKAJTqiSn37vW4QO0bgrstqGXeHk+ujhrmLnCiOb53udA5qxWR1MmHZiL4Ni
nzneRNG8Z88o2YE1dWANYxraMPaf5Y87343U0yCgVwANO2hB7xo2cyCsiKvwj3HaK0YX6kSgHNnB
Hn6wGzAzfwshKSj7J6S8di1CXSEYzlMJ7Cg8FUnWiiOdRerftwz1QFX40gLuaa08yhTU4utdE5+S
6ra8a29454rg18C9342/xW7sWsuLVXwrcBHLbOV9rKZPKGxhzpG6l5ZiutakvhdMpKO2EayVn/Rq
o/ebCM1jg9BSqax7m7OW21ETQpcZvw3FZ+MLsEfL6i+3MF6CRb5jmKMN97IEkhHudt0qTSfZeymc
UPYbpWXLkM8jkY2dN/XcacUqm8aaeRFJ/NnJyOCCPkql6zaWoUNlC/m70MF4Z6z1WEioWS3FXbIU
dqv43FTw6V3jZG9Bn2E9+U2BdNjvOC+fe/iNpBtR+cRhEyBvikTMhpdwOXJ8GH3aScWqCJG7DZ43
VrOq7G3gSZ5ZzcFPDAKVA4djvTASzv8Qh/+fLPA+imztsBX0rZSAu4BH0HVU6/I+g4scOvWSze7v
KLuaAuhXVDp6gExOexmleNueyFcKNp2WxXQMwsylgocgXaL9wsBORsrnwP4lAJAIxjCcyAxTdtV4
PPFgZUKx/DeI9nSu3i5uZG9Es8yTUprateIN/N/53lRBDSnZx+iqifpwVWdyFi1IdO+tL3e5Bqhg
kVYA/s1XaZPzu78lQluqND9/nzwcsUbJuCZBZBgC5N4TCYB8tziRwTzbRgi16hNnwkD78DJtVNiz
9kMmf/c379LFTHwKlDyM8FP2dN4NoLXOYWwUiDipZyGPk2RIWfawLDugD3px1ZG/iqXUcxI2+3Xx
WXiqRsdedTFBOS5Tvs/kNO62rJb5KDdHFtieFuDet9YNf71wnd/Yezrv/CsZJwYofaSC39SxTZGm
Vn//hPJz2UrRgY1RA84Hfs8MAEJ4KLbLh1rKgkXSLQrDt2Q7iHqnJS264/t6H3EI/4lGZbmfNrCX
jl+yMuQfGP8hjI+Q0nhSv3cAaRbYtWrdaQI5gb64r6fLs9ri4PEXhtciu3OfFh9MGB4xZqhGN4mZ
xn6VyU75jZWJBtYqShHIwOLseMBzzWG1ZAU/IZxeK85UyjUXe51M8FVo+yFOF3o28bRRIwmF9AN6
kwzWHaJP6VZTW6C8Tc6SB/x0qxWUKccG+YI0SYarxqB0AD3h3Ji9gBBttR5qFwiCucfcucdNmcjk
4eZB0T+zALAHVcnd4dVvyCSChSAymjHUg1QGKW4yupUVjgCV6TWs78ecZkGhbQEaQdmGIORu3gQW
+gdBgOHWYByEdnxbtwqNNGPBJFZ69tVzAuUyP8Ju+L5Cdgrl0lZk/wwGrx3PWFY+bD0EhsHwE6sG
XKZOgoNFwb4diDtEm7a3FD2TpfcMcbl0r/RzdcLk56EI6IN0c6dJC/4LUg406vUPpiwZqo8lCYA2
OF/3h9xTii4cJla8rzDh7GWsrnv1Lv7I270G1EVRwM/El8P0RFd5FrmKETraYo6H4j5uDcwSIkMc
mJJQZuwm4/E2ieMaWoDtJ9kzB8+jZ7Tr9hsW47iCNjlJhJKDDDCJAT4PqSom0nVZiI0O8iZztV4I
rmNn1RCj6ny5PAuZZGDa6iiXo32igAlNeqCI9D1ku/uA11ocyG9cElXPLEo0AURRmqyFYYxxPcAO
xV+ZrMI7vOP/x43NTbwlQwUC+9mbHlGKWCh2aFTVImjfOlWG6FWwl8ZQ2bGHw0jFhR2vW+Gwmp9+
tuwyLngDO9VFkzZR1S0UrK1yd5mtx00F3SUhKWdMEp+BTLxsWMPJ5YJM/aSz/nk5rDNtdu/ZZP/f
MoioserPbtAog8d7T2NEH98OdKAntxw2Vud9z8Uc+n++SfV6SJxcN4fasjggNiuja9y1Xpx6BZpP
1kE88QyKxxD6fHtyG1uW2aQpy/EiwapjEQU7mdBPZPAoKBMw2gwhlNAo6zqV7ZkXMBrjL6jSRVZh
QTQzLisHgk2EhpfP/vNuILzImqaND2iv6dxPFGxBJcZBTC2yuYzgSsRgCHU8j9mI7C0R7C+DqK1e
d+A2Qeo1BbeVpA2fvUtNrL/LjGx/JLrf9tCxqusnR6G0XITk4MmHTj1FxlFqFev6KfO4n+Z0zeJT
Qdk2Wp4NinoeQaLFFO+5tUD2Qz+qa9ZpbiJH7wLd8UHWswFbwGaLblRidg1PCuifCJSQnZVtfY4P
zPyxf6y5NiS/oiAtoA3yOfnojh0dxF9kWJmHaylu0SvRVI4i5JV5m3oQFAly1+mNuOBYdNtw8PvF
ZJHB9kJXvblGLCTAL+W1zs8t4w7aCyGeRzHgrAdX02gVitj0WtVmc/XZXvF1vp1BzdNOXP8/f4/Q
Tfq9hhMzX6d+r1kT0b4e9KfQLSd7eU2fXpheCUQumVZ2yir5hCET0EvzyhcTBgoWT07c8pZYgLt6
v9wz7m9BoOkVRL3r0l6yfn64QvmKO1APxnstVe39G69HdoNVvI13z+KV3ixg9rVMCuCCg7GDMijk
2Or9/KJgKVxK47ZD23xxnx724/FGZDa0IVs/8Ji8TgGR2McHrDKtBOSJKbzuUV21RyKOFUxy83rT
5CAkX+yH6C12AGey6ntaQ8E4dl73raZw3I6LFxnFEqzJ4NhpE9wKHPzrNhX+r+rAP5TgAqbmQ3Xo
XaS2CameOzHphBCE6a/+dkU9LCvZ5DoKBCz3ED4yn4xkK8WHFTyk/hV6bbCbq9WuNVLTPol3cxNI
YTQobak2Y0djbrY6UcTwPfXQTyuwuXEKLodiTB7pLHDHB3FgQQZlwqZL9FSxFWx5XpTVLwhUtes8
/SRlrOIXem0ftiEbgVzw21DG0GHWIcdzwdpy2SjaxjmZGK0JK5gVhRv/G+nr8WIt2NQCOcTb6BS7
3SjvCoS8mhMw/CVv2bK1VGDXlS6KnSdXvJjBtRm2izZQSKjsZHwy6fi9TEn1IJMRdYToeR47jVVN
pVFhEmuJ4MMfsgTuvmkdwFYSZJ7eUI9egn4LiqeCCmqIL3OO4HP0Z46ZFxsrqE/ublmEkkM05q3t
oeUEXQLcAj71WQZbp1MXf9/xn9yLpC44NyYPyqiJHjrEH27LRpE/DVkOUouWwe8tmXtD0950Vh3M
F+Q68uew/8J2QuCGDHdBpjoB8Dxls6DuYH6bWX3AVdLkyFA5BJ667ofu1At0MdO1lIvu+0IfpW7i
bchUBaIDMLiIkr7sh2fz/XYFfhjSxZBAEfURjb6PRia+fP+H9WQXGWDHvQTGPjEzK6oEhSCM1uvT
y/WSM4qdqoOoAnfpyqZrx7GAIE+OEFo43aLzbD5VqUwzJ4HDJJxt5IfUinvZzSc/lSLAlhwLXLxe
ANfo8bhcanxNusgku6gmJqJZpnDK11RlrGkSIeQw8UyT0ozSnM5xl/kWTczrCJsEjc+yiBEOXSeM
xIBttfpKov9U2PBoQkfQ/YnQqQGQ+d43j4LKss9oW5NeYd8H9UEDzC1pI6OEliH85mdDZaaH42ps
U1XFwqzyhtuLCnoAnjzQ9XrRmUv9Ol0ZGzE2Y/DvbwX7fnOqYxvZrXv3pHKxujRESW/IRfPfbfA8
786kX6SZMmLCBgb2bV2HRxOxnnb+fcUwyhFMppe3TBNjWNKBetFFBrw1bxuJfkgyou73UgrnGehB
ayyFRmj14osafedvpUcFNFnFm1ftWzhMvijpyof+oJfbK9ucOnGoEOqkcGRtjSJZZwtfp4KvSJeT
NusKXdHTl7c7tLE7zlWqnMxo2Fazu7DdPAaYd9jPsB528/TbJz2SxDJLUyInSFIwCljNBVso4kzW
l1DNJJcBeRpNo5mBVnivjZwucZHPmJ7c+yTSGBUY20fRap/HKGtIt76JqpLNtS160WxpZ0DvzG3B
W/m+qrwC/J6aRv8MlV5f2K9ES0/y+RlgU0LHJtfkcJdFpcNv0O3UaaDgncwEMazJzyFVkuL8reXI
nagzQp0MVKQlQ8V75k2Ji8DNZYr1pn5uxtUCr5oWE81z5gvuqza+ZARVvQ96ZTPnM9PWX5SIKv9R
DYzjHYjxeNO+CYA35IZjO+J4QCGHkZMHkNbLXJT1ThQELqdqqb9xfCNNReEQV9TkEh2tlWT4Colo
Avq9SqyH4k2xAdI10YNnY45yfzeRIgPKnU/qIJXdIjsJbTXQJlm8mWdIfjKknEgVIJfxDd7fC46e
R7vRQWB14u0SqWMv8c97Ylhxm2OsGDejK30Zud/xM/vLliOFbJJXFjFmxxF0cQHsM520rpJ2bRq5
D4wpO6ePaeF6GzjaI1oRYorlv1XK0xqIVsJmnrDIHGUN+yr+JCQVS1ZdgMEA075kULmXSlkAMs5H
tmFGjnD53Q4Z/NJ8Z+r8G5/g1mlOqtxJamXaspgMDfE0uuml/LUyik/I77nxx7hZX5bv4PIdI/Xe
BdmEJb9HKcSWgEoWXFt734dA/oMWJ0c/DlGvKxzvix4NlcdUuBoOIsT+7YOstUqIAekEMBf66i6n
Ng4R4hlufbLcUIdWENMKFQnQLVQM2J8TVroUGYG+nnD0aBHyakDPaXNV3OnchO+nNLmdywEaxzib
CGGDvCZs/FkrvKa8Kgz7ZYgrL2+l2je78ZiJpxKFDu8k9mIh/FTfZgjr177xWXZSxCbRHrVO5toa
eu/OyGG/d7LnbNFFEcQ6hIwYjRkPqV1Y7e0acIXBP40VGTrqPkn/mmcjhk9RRgW39DFbBBeO2E8P
Pr2BRWjithhknns6mzi2jzmt4w/3+jGny81florFNeLuGqbyGp5cxK/RKaX4T3LBqFGJSKY4OA+0
wtMuCt627Y6/9AIkOCH8sHCLZ9RJuYpmh20dIoXRJXxpUBd6R7CZWYNEyMrpIJerLn7X4M2kBzZo
yVURzOaHPSoBPVrOo/a95TcpGAwL2XUkLGDEcdLUd5WE0CrdG+5Yt7EHtvKBtTLcYikf0u9zLXtC
yo7b0G0pS63G7nafob8ZOFEf79/RrrukLPq0tHBI1bz3sbb+3BCN2q52uYObcjrIJHZboZKGGBII
ToHWLahuw1pVHa+VUk4B1OELqQ9tbxdNEUM/DXRROfQLTsH2cmzxN7guL5PLmsJzQEpVhQG6qadJ
aj+wibcf2eQ9uLWHF6zGcz4re2FjfiFtoXa/2lgxbm4wl9M/UI6H31tJS2Yy7E/uh5PY72Rtlt3i
O9HquoUcIWTDtSnho4SXt9X3ROjY+akF1GYPzZPgW+Hbfiqh9YjhdND+q5xoTP7X68cgzRwQ/TO7
VKXqN2jUG8MWRsUAfQDqiv6Am60mdI+OHavWJbF/haZLvb6jxpADWwQupM+y5uuuyhtNDvlkUFgk
wlv854wF562xPRz7qQKMVL6+TfuSjm2ZTZPAAqBwhWVAD95S6F7I6HCGlErHjNEDMJp4sUHJ9UhI
tJMYzvaxQptIGpfqnw4DpVsfvi/FaSj5D+OlFge3rvscETULV5RUPbCVIqGYaRgT8P8l3naxQ4n7
xv92NtPIkqfQo/OQTqklUm7qkUFObLvlg4bz1ZgDZU80LXNtisusJXvafRE3DgUAsNfJgpLJdZbr
dxpXtno3B4XUWjc2ljcunZLBVgJPZs5Z9UtAcygoL3iJqezAzl7KAo89kwhuLwrnlxp+aZ61+yYh
Rz0KQpd7Vx6E3q1oMicjpARgdAcIcMDZ8ophpaLnXwZVdP0OWnaT6EQsZ5q4EzKatPbG4ifcuoY/
spGfc1xakUdDcM6tZkDg1i97MVdapN/B+CrV7eOPBOVCYGl1vxUssW4enXFDK38SIBkDrhgYe3Sd
XN2oz72+OYYrL5bCSY+Ws1A/sUw359fwa2GcaBwLONyXcwPF9O5G9E6J8jZuPgwazMKvpiJFS5eB
ap5bURlb9e72nQ2PtVuCNUcgVgQvPvt3O+dm09lZr+OU2MtVmTfz7mMpDbe1fCNp6ZM9F4LffqYU
Ls+KA01kJeB2y9YgI0VfdAqYfImKpV1cI7zr4X+nqmhPSSX35lKHPfnGDd1kkB6WfW9NqQ1lGV7W
jHJFkroRCVSyRvqsIet5Z0hTSPJyHafbAauVaERf5ysyV1v3TX6PF+T+Bf+/MUbzaSGaxx+vvMcV
zOIst5gQTb7kajckwbV903EbkrDw1OcknhkAfZ4/cA2hnFxaL8OX65eeuziK8u3LjA+p4Xzdxc/w
zkrwuxWdR80NtErOniw0y5J8lxQyWtkFJ8FnWG6CclmJ87RxNx09wZGSPDuW5N2KCF6eMiC4qIIp
2BBWzbEFFLYw7JNqG5KViy/MHveu+f7iFn0W/aoZX7uJ0uEbqacz1dv+Q/OvUMgQpGvDmYWUo1dR
XCCIWsW07wDNprGkD2BnR8329Z4gNCxdbmQlfaLfl8ROjcZ0FxvHF0CE9eNRN+/2wYNKP4vdWBan
J3PiY1oGGBDAq5wEIuXa2e9BYizVSSVlIyYjAkbqebKsoLTk5M6tpGftMnmpNbQXRNSow9AZ+xhH
EzKu9tbojgtgiXw9my+NbBvW8ACbNlZe+GoC0lVCpRK+sTM6J0VAzvsAxGKbkB9mpuLKZgNd4nbW
kVrI3qEw3mNYiuHnAH+GWIikZVCDvCS6yab/GhOGwNCpapxmsCdFJ7rihWFEcbHh3Ve+qgVkBW2m
dBeIqUwFLKx7QdDm+sV00ERFpO8AdREhRt/FZiAfV6OSyI8htd1Re1fqeCPFmpUR4G5IiNyQFjAb
GZ3jQS3gVfhMQPk5MWtn26RX9Y5yL18ifERAYodehXCkJyw8IvMjs/Np/xI3ukKTySGrOqLMcxau
7NRTZbHvkEdPjBwCDyub+P7UsPdrMVRr0z5YoOyAoavgnhfqATLziOZjydSnvT5ym/7qYzjNtBJz
VQQvVcFoP4W3NIl3jAIy21BdWHDkOpw7G+MiBTfA/gZl9+8A/vY4ckRlPVlP8cZzvaE8edWllLA4
Q7ojrgr1emuc3/c/P5qZKlDJVAy0drhhc4VOtwi0WVMW5kF5mgHP13kn0opoJVRhHFp86K36FvUV
kEA9GcwQsIxP7b+4HerrYR3W/+beDJnj2fXZ8usU0lMuNuhIOJOdNzckvIudRAftKzMp5Tb9pc0g
A6vyMb9GR4N9elLboRxwwkTliUQ1o4fEeF4XFAzlDbJ4x6b8oa8z9w3Pg+f3IhBj2fe6lbv61rX6
r7xtoNXMplku/A4Z65WUxclVr47SOER0mzvxBLyW0h8pxk0MCiyuC32xTjDBC3sI4a2fX6hJIhNf
mroJTTqXuV1BEE71HbVxFd1gPVUdi3xLEyBYSs59yc08fQyE5fr9GgrEDvhzkHv5dwiJ4wTeNEOr
FVDGx1mA8mP6Mgtq5E3+zelExLEWm1gm9bjBrYkc4eJ6lae+YDjokQ413bH23pCJK3JZ3AeGk9qi
21sotZcQYZiTPV6ti/wpEajSWDQmCEdNT+h+Ya4cS63V2zf9aerrP66iPw0/dR28JCRfv0fqetVJ
xO+dCrsq39uKQAQekB9OWVdFt7Y0pqfnG/sGZ2X1NLScy4aXu2Mn7GJ8udVoJU2kdIsU9e5CZcTd
0kBg5yPq9d4KAdpJ1o1OQYgJZ+/oD9ThbETMhVFrQgd9QmRy5Sbb6SrofYF3F2urqWkEZzizWmtd
8TwauKhFr9B0FC45w90GCpuKCxGLNZj6suMMpck6G3ee4g/u0HRvaViB68vbjJzGsnv+hxx4uIo8
sxM8cbEF9aBJrArY8N8bWm6xD4gNoM9zLWJ/vBbrYRxHzWGvuimwEpNIJ7ePFNLvEmsZZyo6ufvb
85bI07+BB28Upa6g5C73ab79JB7wdyCMXFpq/0kDQUfL/fJmdBaYDnAojngrTqMMxApUpmc1fLZM
UKpGyIm7XGXiDrADYROlJ87KKAIWP8pbkP6O1vOD/pRBq7LNZe1fXdHoUSn90SVAuVoZ99RlwEGK
3FoS5icQC9gg/Uj0vGpr1M1B4vS3zAWRPY6AXfb86U946Cm0BygtH2p/EE1M4SI5Qom2wbZGzSpT
lqTykLWV8oWZxjOZiKp0IDfD2BFNKivU1vFwyZF7MRiArxuBXKj/6Hdfie48RH2S1n9hpTc8LmwP
3bRlgCMpeI/U1ykBHEMK5WoC0SF80gyYffp50D2I2uJz2OShMPvecvs2zKsqcsgns1W6mh4PPfAp
6I+XMFHZUPGoj8w3V6h9DeeTHOEObXkkHw111sX+8+GvvDIbXMG8M9zf9qLefMue+UO+PdRY7lXJ
vqD6injGbwUkTa4m1isLxRl+zSRviqFh7infFTLrlW4z5qJuSr/BKLg2JLeVUuEkX0dm+yeGSneZ
dtW3LkS5zV/kaqMNvbxZJp6oLfs/FbVBwyyQecrR9ahPfPTnW5qFVBF3sHvJ+r4EHaBs0Qn+37vf
L0xhVgsd0tEVlPdPZ2y529IDa4z49MXINJb/v5qBvBgTM0Y19OwWDoFRQHEqWCkCcOJiIhVYC9m/
kGlpPhy+JJeE92Dy0Hlg9EIqIcTyuuG5jVeTFB0vaaAPNLuQkIu6lBkAyH3yGcMAmn4yvhfCvS3F
OL1ie1i/nPfckGkvsIYRNIEYknmf/7prRBi3vGaHTf9FgejoQ7OnvON7YMJQbW/YZmzF329kgX47
TY1HMAfakAIazuoY82o4w9bWqVZUlMHRd1qbFKEyEu9n0k/qcXiG7TkXS3yuyLISJCjQoe5NwTfR
lChiVC2Sdz7SzKhpN0MarBQk8CqPWnnoFUKi663s5OiIX4ervmoLNAVhY8ZBwTgXTl7NtZKmZiKp
/adTNMIaaOZM3g4crqMzwEr3IkpejH+RkL1KmblqTQJB+ulSe7C5/fd3/bjepuFKR9s5rL4moaQo
65HD39qlNWaLaY50p3RJ0FuOKY3RthVGofcLMChL5dlaKj7tihXhmSePqYyw/2hsW3KB2+lL5DXJ
dZaDAOsgyeCEmRPbCPnGfCXrdCl26nFI6BDYGLQ5eX6rhFEt0EFLq+cEmzb35AHdBT4y7pwc5LbY
HJ0rT+0ekwK40QdSzEXD8qhWB9Kc2u0WrOQxZM5NzUD5INTe80TRVm42itlhFKj6nuE1I9vUjY13
6LMw9bv++2N6Qa+vBfGk7g4eoW65K+8mmuZpA31AE1zDHWZq9pg/wsF2hBYUANioN9A2KopoHn5I
M3/NZvnTrnrIr2BYSzX4Tvc3BzJjwZanklV3LfBlmSjTzL+Ff6f1orw3KitTN/t4Tka2R525in8B
ojo86f/aUKbm2FS76fqzKFuaeimI3L0P6O53b2zflLAw1qZ0fBRnuKEjn0+XRK6CeJyfwzjcWqe4
e6UHep4fAN7vUUw7kmmrUS3Rjav5K2QiZo81u35MiAS5NYbKdvm8Yj71wFjcJbijjc1INVHJKoJm
6vk+fKlP1FnnFgLM+w6vg5+dBW0gNT7CSOY+ClWC5hmv2j2Myj/WNeIxo8MtbI/iWymo5eQ0Slvz
5PY4n5Xjnw83a2jOO2vWhco1ubxwYjKONSmpypecqoEj8DIsjzJSwNmOkR+5/gmRUOS2IlLhOgqA
HxiwWFzmnn6PlpeD+CURt+f+rtwLP4EILHFjA7Ig+j+G8I/TK1OEt8FIrCXSZXWfPmYHZmehfUCJ
22wTQOGbXbP0LziTIIKcGXcOipRuwqFvIq8GLc1w6f3YkX20XGcmzVegnyVDQMJyhqsAKTCD20/A
bouch0rVGEpjmjtjDCkztEdRRRsY2oJGN45D/TmbQTsnz+jeLNlQDWCeczlSnbT3iPDeKEIJfwX3
EDlqLGTZK7Dcm4a+NYW04kYS0jGSEDEFJBTF+dgpS/16GTMmjJAN5SOf/egq8hhoL8AeKCiJDD/l
nxXeDll7o3l4DRWxqzhzCRU+boA0G1+SqhJehpEmKIZZsOKvLksLH0kvsh7a8yRxWcQDj9SteJou
6VEXYwwDvFDPD1buxy4d1t17rtsRMlUJmYKU+tdGcu7ASU1EJ827zZ0/nHeDtjAcJFYW4zM/BAnC
1zkOGrioqTba5YRg/0/IiIsoBlOgPjDNIXA+aZPnqTcuuXIYjdMP1ZErba5SRunRhqnzcoisNBcI
6O4b0GE4cHz6BUvbWK2Znb1MDBcUVJ4lyNaPz9ened7HpFGeVCtySKYKoN9rij6t90R0OSYtZpdJ
03N+RPapRzPl8yqzmjPVCqQfJtLDCoFP96r3bqdQbQDmQaZO4fQmH1gYvQd/8YHIzWZpgd8c79Pv
8sTmg6wqOBUtDF2cPxAA83qzIMwZ3zAoQn436ajhloIFWceBjaOWI3Gt5erQybw3wAwFaCSl1zSQ
nBNNXVxzUmhiuO4uIsv7Ei/AyjMu7k+bHPmrmO1XNUIHD4Te0a+Dv2Bgs+yk6j/PqDoKQM8TGSyb
4tw5s2VkzUghqPnL+wgNyUApg3QouUQ1ROcJE3gGW3ik5vyFolDbQcxoORrmQTKwkrrIM99LgT1l
aYFYznIhOp3HzcVvOziP7p48T6dRCleQSf0ZwPWQWHHUhQdfYyETXDNNtOKs1KiqK0V+kM27XvA4
fUJIcxNngyxtC5SG8ivP1FzZLyZHrUD+zb035YqdIrXT2x0b1iIBrZZbaXAEER8iWeZ0/OXoPVgC
AoD12ScMN/rgM3koLsN30ZBWfFr/MghO/ZhOYY1pe1YcuO1rCnuiLFHpRmhdLvQoWpdFYSTER7Mg
WAo/cH2zyfUFc/vi3DI/G4kiplYUatEk9CMdTOrOthx5MAtoX7oAoG8wRyQdF8p6ip6atgAmeTji
8iL5IssU1Q4qbJR555fCkSW0I0TRuWx2sTjc0Vt5+KLZ6OmdLFeARyBjfXRYTB/nKcqp0zJlgDvy
RAXJWKuj/hBV+yrblTl6UkgRKgEIbrJ8sOieWN8t1k1QcZRMFTANqiyWchNCyvK7vOvQXImbr2kC
LIkJsW70S2LlvPtnAEWGOAe2LLkTARK/Jyz429e2Dqdyl/ZgAGUm/w9y5DOX+YvIGnaXYUAQ1BkM
jmz54u0krE8miDsAcGPep4GW7y4LjBUoG2Z3YYmWXpZtcg22X/vIsyWpeaDUUUYO4uK9iaxPsFi2
EPanWEHVLHgzRqiD9/5GHqWE6PUR4ThqNIHamcYBMOCADNDHpAfanr2H2X0dbZeHPv8ONK3WOBec
PuuEby97UusFV06+ujs9rgOgMmgbBo5u62fyv9mcsLKNOlSccrsY2HagU7T6eQTvpmr9kvhtJV1J
aqms0D0pLi9D37zF3hctsAwgz/t87afMfI43LapnNfCQHK4SKYxKi4Wsn/NJlHfT0bxuJnAWkgz0
gsT++y6LPTRwVp0HKFPPLcSZxsXRW9hAaCWI/huv5Ue+YJQ0cV7TjgOwTaJyzDwe0s/VX1V9irll
K+GXtk1Em9hh2p3kwR5eXmSCJs6+bFQupbk66KzngbrPlHGoqSvpYs7DVRR7ED/BzrIG6Ur2TBtT
O8LJSSjFNQY6pyyiyI87d2tH3MJNhm3RQf3tMup5gM3wQx6H5uRKYk0MWLKeysiXm7qZmGBQ/wYC
1XnjYzPVlJwMIDseVUEL/yefsJLsTfSfLcf9KeV5L0wMrNHUXr1c+zemzFCWpyxRvA3RrDE1Qd1v
DJpyj61Zag+BoCFERFGHUTya9t9HVTtxZ6YecLpSR5xNkMSR2mlG/c/oYM4hq3rL7Zkdhwu/myJ3
yeWk2mE/z8t6rLWaX5IhlWeWqnxuWXxoT0DP164O34w1uCxWT7M5C6DaLg3hXkpTUV8MOHnQCuuG
g0in2ZKyL3izV/GGyKd4Mq3dypWu8HJkThbyn+sOTVpMTCun6JcOTvPZ0nKIZ4yNsZVlAtoceRR6
djwvJBYl0zeRFv01KQ5/tuVuFJaJx0Rvupn7lSRq5rsiNvE70/iqdBqiwQLzriEP8EdhyTRn40Q+
u17wTYJpqGzu0Qvkomj6sLKonNaB41UwXjy20LmmKE58ZzXdvoIfwyxZ11Mjt6yBXgr2NoH7mbu7
0PXNRYTWcgHIRBf+w6T1Qev1/bOg2HxtC2iS638PY2jeaL21yWM1Mq+TGOHyBrJfEfSfjd+E4ZIr
x6oUClaI2fioPc6ZkKzWRj+sil6BnARSYDQCQaj4weSdPelOfXNy6iZVR72Q5v0ga925r2UM9f/P
79gKa4VyPn87phLSliXSkUPGOKlcCYEsPYqayaE6K5inYCdbRCYu3P9Itt67OFpMBS1IGiX5vehv
1tu8fcuSI3F55NwJnGA9OaSW38ptCwdIL84tNQVeFiFy1ZOh9WQj642M7fPWWKufebeoUjhfijg4
XLpzoAFLHNhSIbNHbA2YsnN2aJfSiudEy7LgfNdbMfU8rA/c7ZgkooZaxbj+5uER97s8ibQfHv0a
zifFJh5e8LlPsHufD/rgak8wECvGjqIqfiV5KD02Nyd95LXWnlFqo6ryOdZBS3gY0za1VylS+E5D
pcgnt61tFzbVAtkiOJseMLzJrKfpxP5NCVy3qwxBcJSIpKURt0Mj5EPwh20wjfEnCxyph4dl4IKO
/GKJG4XMM/r3IM72nPCa9nBOG22kBB36/m9+SD1h1FWDaXh1xJQn3AXwJMcppmz2EyeK+SruSCJy
dIkcpGzv914ZZKY8AfwvbU9GUOrEV7RI1bx4tXD725E7pzl4rTXkj6db2OK4ZXpcVuH7az0GAESL
itB7Utn5AFK5qqtOtp9izQBtOGSijuxf1rAgMU4zjsJKl9m+PhQccjXsCVe8t74nvqRCDMaf4uSm
8aK9U4QoKo3HrkXGtdix5Rma18GcKA7em/F7AFs7zqoUNPmRT2kJvrVpDlcPlYWDOa7yMHGtcUaY
kq0tXVGXRw3rffCJpI3ljvKATP4dAd4M9VpA3yAAMAKRKQMPMiB+iAS+EX/Oh67uGZ5e1n19QEkZ
rFbrVmajvSXsMybxRu3wW4zKIteRsrAs79lnBrfy8I4Aje/jVlOm6QKcW3etw3+5PRQ0+mznMm78
ZsEzRe27NjcEapnaOF2JcWNdfGH3QZaohNJCxZA2kbz9M205ANu4jKZ/9VT46NQFAhD6eqk6Ckg0
jt0vVRGjJMB9kXrh6mR3XCPQiF1ti9W91YO/XzAhW1lmpqVg5AgCz9aVmS5XhmIW+z4XzJm0DT7W
ZKifiygevElOheyEWqoZj8cMX3WMdcA/i1MGuNAClKdgo/mJAnGn2jXSQ3fI/gpeliW58HH9z059
vr2e4amTX67wtMuezupVscbuyUKjxgG47a5RVuMZzVTyxG9YORsW94qvVmuShT0eDYSILkZYxHcN
w+ZRB/nh4611BMh7hTYElazTjMismBSLl61lYePSJ9/IoTg3p1uKo8rH9DBNknGOEvFmRqR+l6vg
w1aQSjAw5uj4Tr/YkrH3QZX4ILuPSP7IvpT3DT9PyU/KnClAaIQuyHMwJrhYgSEPc4SpjdCSLG+g
yMfOpEu0y5HGztcJh1K6XJQZO+KNpR/qwouUGVjAzWG13WP8LuNBml9nh2pmV4S6rkaGn4LT3myo
NK8UX2OLnIt2tXT72ufFq6m19PlY6shAGWtq7rwUpTYy1T0njHoVst06W8sV9lykthozhStiS0dB
JJcxXlfpSU6OxHDLSI0PkuFXQ5QvivlyyvHSvIqtWSIEAuTm2LGbcXn8Ht0YDbbDZhvYisejF/7W
e/MV1qrtvM/ptIze/YPpU53Ouz5OUJDQV9tULh1h8vnuXDtlx5UOfJUv6Sz7Mk04VPalryhJRycj
uQu/uefpaR7jbh3Q36EE0J4zTzF92KSZSBy7SLc3YIvc4s07FEtRFV7Y1J2UxflCqzTVL2Bo+9Qs
qMju88YwYd2r7YMvUmB5yC45L7F6U03W3YmbWorbBM5hoMznGOfIFThOXXdKDbgb9i2VlqHG6HY2
psz64C70iNKlVxwHqSqtGkE8YBXaFPiHg8qZA0AsTKTFHBmG5xvaLuSGRrCIuNR4Ls5RCyjytCan
32G1/uKl53aPEsP2eLMoObx4FSssnazGy3fn3F4ZozAKIqfq7Ir6s9JgGRsKZUI4KhHNlgjzesOu
OWlXFcoS30/u5m1hZeLAFbsMXMgISXDuzTyIvm1lW0mBcvkyrz6HveikGA9iAJTMEC5nWdw5RiC6
Ef2Cv+ChUmTFlhTRsekclVm6w/jxuj9WjNMhwUzJifT3ZYUmSCjzsSYd8du9O6ImAhAAhaNeOPvN
Nim4Yw2THroo/Au19Pq/198Mj5of5D80K4xjA4hIH/Uti6rZtgDjfILzLKllxvAzFIts0pQWceO5
xPWXu4zPPQuonxwNtgKvhdL5vFHVhYT4e1f5gyX5bcCcj6utC1gpPI8Oqg+e7BApr+XH6DCMYeEu
qsVCUaYvh5RSheubZ1jOxEb5jYVL90tjS98C3+5ZlIBWT2Z53lNa3eB1h9+fxs+ClqhjpLGBZbCj
rmaWTtzp7YuIJmA6KGL3Rj3783EWDtA2rORSTpJqnWN8prwoF0+6aI2IBdEVHNL+f8Cx4xzHEpsK
Ha68/8tVNhnIXGOI67+0UdaYjoT5ZBBK042RNx/Hm5Ljy8EfcMPI5j0dRv2DrGTFIxKTVyoGOx6y
aw/ZnGW9WrJmkmjvVTbctBLeWueLZZDpQA1V3iLoMshVlu790pNZ7xBYLQU/bKzmArcQ0xBsUWuS
tqY7e738Gsq1QJMS7UecLIh6zDoUEZxcrINNL98S2AuFm75iWrBnBNvjG6zkftmurznbBTFTZaia
cN86+M6tOPiKaW6QAR5YJ2DvKnRhzYBXgTztnt3fNvNzd/IyZ25Dp13sU/5Znnj0BZD32yUCUCkn
fIpCUZgLZMlMqEtauuDJyd6ZCuOwEEdkJ8sP+FwBRturow80iQ54P6eSjoiLfPOd18rGCqZFoaVs
Tb4ogArrGDwN+WJesWPYtoyvR8Wjs4GqZTIOIYms++GCQT1C8JcjogBycCwfJV9OuopWm1kwwNQW
dMIGFEeWSiUZvbZ25atlS34TcaVg70mTsJGCSzBKzaiHx9N95GqZO5xyG9ZDnspyTKeV41DEg767
ui4PtC3Xj80VwFI9GuUNDlirWV/XdfxcSyl8wgoN25y34/3c55U2YY/ZL3ruIqWvExbiUljfcpL2
3efLMHQbfZTM97quJFTXBrmHfXHhwCoowhAr6WRd/uCl7RcKjn8mV7w8CAOd9Cp1edZS79BI087b
VJVhDsGQeNuO7CjfBO3EAOP1gdB1YkwOq7Aj3F0l5ohiPFPV6ZHUH1TZCRBw+H/EdWgFLhIDBj97
wP0Gwfi/3rjwW23zivrtnttHbo0yVxWm9kyqtMuKCtxeHWN2Nm4E719Vg8QTb4fGmps0N9GHOUhu
7CTDAB3DJof7we020AoVJW0JJWlTSpILXq6zAJNJOkuyFFHQkSKWWmyO6jmnt/kvbhIbObNaCJGh
c/3LIu97IkcNbVFsPCjxt3qJgWqTW8r2oIuTIwYtgzq2lfmeYqS5HsGIcUre/+CjV+3wMlBSDs+s
4KZ5CiMbVDB5gVMEvgQ6K8tAareJdEeSGtQMwsRflbx+tbxGB8fZ1Or2kb4FRJKEtWY/RrMb/gYH
VvVBjBAO9RoqIN0EK2UcoAJqj699TUf1TRdx8IUUo2ygU46jKMPyaZjeiwEC1oseeIr9xftbvb6Z
T+QkVYAEgFHs/1sIXBW15XcQr535e3ae3QzGW4XdKGkWBpBM24WBS+DgqpginVqO8qiLUq6ykLNN
oO7X+4kYjNwkzdixp++Dv4oXrfUEE/PE8DJKya00KciJmJKDiu0omNZJoBitXdu33a4+sEx55vdW
GFN1S75f1IEMu9rvWJaTSg823Ve2AbBlbLIrclJF4DFdJUzbXv5VaMqKkcXDfgjb+FadqOlbZ8Ye
XVOrYY4L7+mr+Hcdr8iqvp1SJ/RRSyyhH9J4DsBKyNfZ0G/Ba04dQ7+55Njd78NX+HgiIA6BZ+i9
Hj60TO+UVee+zgPEjqukgsmVCIn5T15Znw5ddLKkVA+Dnfj4c+OqyYeUrFmrWa4Bhuu+J1q84vYV
FrjRgTCLsBIQHXSmkkIh8MU2Ct2EEcozMXnhLGd9v0kzhlFguxHAz2b1LqWcTmNjPIozho+EJGhK
mD4C/4cvAsbywrPZ4FsA0A4SsHWbN8zjImnSkwP0HowViR8PZUfVx+YVU/W8i8fV1IGMWANTP5aW
quI8IU8nl/cQzpLpP6OZHMjbsYWAtBmSVyxniES5p1FKi4fCJbTiV409kuMLD1Fr+ezy+4grvjq7
XdxqKGXGex+Je/2xdLY5Z1FJTHK7e9xdtxjQcV67E7KmcXmWacXUtGVe6oQx0wOAG24Fan7ivK0c
dYrHxn7OP+AALCm/khl6kDjLGDeX3liYTwU9O+oDKjCMa8TQqJHAhgdyXiaEQkOjd2MmmtaykAlm
VsPoLRCabFIuGokbleu3exSr0rExlS/X1FImEpMAy9gDIlk/qXwM+n3pm9HGQhH9QEOgNbD0a/jA
HDOcVPv/bqBQcRvd1lei3pQupcK76G9K0pg+uVXxOgaIUQ5AhEUNIfhhpxY+gL8zKNzNPJkDt1/a
Bx1scpXszdRHmsPg/NGJnC4DKhSzfv2dFuFVN/r8zKF+4l25WEWy3psxi3h7pR5KaN14mIYGvdvp
vYrXw5vrKvLx6tejzO5tT8qT4Ksf85/bC4qmGzrx9c31+mvQa3WJCKidX2rxS6AczA2V5Cc0Cu7Y
4mWaAyOYVP9sARRy3smDEeXVGwMVX0rsHj8/UhJa5u5lQYFSPYtWTiJ3f/N0tDPmuM2iDqqtm+SY
ufNReDU261jxK0gM5MtOr9vNvqNlRldusChYHoO+2Dbt8S48jcOw+9mdK6eU7av9juem1+x3yhyj
7PPLHroe1XNlNTKhyL3jg9JhNMnJt/Jg5tW72JlxcEQMPdeKuoheYf8UTB8RJ2gUhkih6sPO9DH4
MIDC+ZRgSUSo5uS/04ZWaxCUUYru7zroKAbIE87+32hskuuowKuMwgvHIFA80DC0QrDoPl07fyHv
Nc5btAg7HUL9gTRRupiMCmkcc1iitXxPmj3BCWFMgXv2uJh7PpJzA0RZY81BfzwXIbHZUuZidFHo
u7il5zH/+lPyTgbkdqdynNRdy/B1YOm11aKCd3CCyG9mWpQHhg8/KrCrvot8GGMjHGNwxE0UHdP9
ElTmk94LEkodbIkxERrvhfOUhiLX5gJlByS0SbfmChNNqMofyDkuxhhuX8QdIvgylP13cdpnpFAf
gUVyk3dKt87QgTWVBPjvPADXzqEK1rMAR5zSwNTeBK2c2d11wwIhjOb72sb5WD+uMtdHL3JUmEPX
A24isMWU7vKD9eZb0HC9Vpt4AoDuLB8XYJlJ7QA+Bl5suy7RoPI57tXTNzzT5W9gAZ3uZoYtWmfZ
j13SzfruMk8JD+BKHgjqASDa9Im0LaNqMdcnX/mugzWkKVjRySL0Nxqu4Nch9g3ZAc2sdG5uzgZg
Y1QIozeXsg7TwJ08uFcW9VGUqv4188vOmi5piWIiGHQ5kVP6hJFZZQuqIuJEpwkLxw+p3QZXLIc5
9qnyyfyUfEon7F9WH7tbf1M4Mnc9O/f07uEb/PWRYSUe3ylxswLUDa+VCtHh4z0+br9MNztTisBP
GXblE17tB0gdy5H71HiaOEXl4n0/Y3x6B5urG+IW2oNoChsZ/nlotA8xxLpE6O6Dk6a+JoxIDLX6
wqt7AjALIke1L0VGiFE1HuOfCXw+QWD3n4gUQsEXRf6g8/oGBI8uX7136DbydVXifij8BWpmIXG/
B7pq6hxSQhwkd+nzE0WsMEGWpzZcBF7/Px5vm4hB7ZmZGirOi4nZNZMqa9KY4NWg1w3t8Wyvj4zP
ZO6rq7Y6AbS0QbfNkL1IVkRrVZxcfAdRfI95elaI/3Wkpq6jq2fQ5JRuWrwxLPx43mV0BwhfmiaP
bEOdVZzrisxEPFI0lDsaRZj3WrKjI+3P9BZ7VZHsCjCO5El55uJ4DmVXADiQ+1AN6QqUubEmXdQs
iR1h4LJvhksWlt7NZDWhj7BOWkeEPvBrSwrzHlbtKEHB7PxQcZ078CJbcSbr3LN/TNBV6hlsENlL
7Km6XQfyY1g0A+t/XUVL+2egMHsr+9asjGZpMiiwvLy4lBpt4hPtQb7Y902vn4Ni4vp4310m49On
FONiuLnptSW7/WjRhdi3FkJFmbRo1hFOpO54F7OmdwqyHSNgAfxkFplam8bBIc2ywrXRgQ233WOa
Y/dmavODRtTdek4uaJU//RmTW/eEm82Lux8W5z3O4tNfXQRK7M/Bx0mYGmX1RS6KWp85ooCUGMm0
bZOj5XmuqpP+ACCppnO5p5SWXOWZD+VbiqZxRLCL+CDrq7e5uHWCFJ7zcXwhLoTpO7fNRBCp/sL2
c+2we6COMLlpxBX8ABpOmabxgLhb3Pp1YyZFAxziSz/VIyybFMM+FgOD4qYdX2QLQLTfg6zMheeF
yBuWuMlolk2xtpT4p5UFZiWpXpSSLhWOD/mLOiD8pNCERooV6M3/TNXZQMOiqCUKdJ7DPKGPIdl3
UyWXQEBoSH3GUGFEeRGoB/DromDfZNsYpeSdaXyadYQ9bgzAIV2W/2u/t9QuCLENcJBIVd7Dwk0G
QnvI2NQfGi8YR3F4WxQ8iPzv7Oem5OmhyfMGPG7+p3kL9lzXFeKx9BMhueL1Rql3O42J83W4UoSN
arBr6NPymIxG6f94n94pN8ngX+85J0tTE6fVzbxg2M/nruq3abgADCyR/TS0E/48rfHOBjChwjXX
nLv3BvyACNlw0MKSahu+pSByQAovtAlZO76VK3n0xxcvqNT4cTwftEYrN54tmph8HgnEEgXTwsuz
DXuhDbJvr0NJbg+BNscRVI+9zxFv+fAHVcxTUCfuZtj0nKmtXEvMAn0GGGpJz0NStirE4w7K4xmU
7NhSnFruPAktC5NDdmvrTbO6mihb8NQ2d/FjVuBUcTV+OkKpvJlZoCNuH5Z7fysTtHMmHILOQjCz
LbUMQi2GFyXKo9x1oDDGpgklT/DOUssHm8Y0HCKNsVG8VafX7cR4v/Tutz7e2geMzeRg4aJz3Prz
xjgTZZNYK4P8sY0SohtlRqFrYz65DaBBccfHBq84uvYiuFArQy8rEha8fHCi/Uv4LW4M8tuVoZfg
UMSSpHQrrYA4fWxKF0LQhla9qkP3wOgR6jGfXKXZQjyxJYWU3FblJ6V55fJYO2oj7wX4NCixwvLT
Zvds7AQIRrmvTbvkW76PTCzxaR/fr9OLAfgLVxAHeh1dkPwwVc+mg9dluA9QjjsKkT+gU9e48kgu
iBifjqKOLZHKhYr8Hv9DoTvVlO1V/JYVcI3J3ndY101JwISj//e59+uc5/+zeDYkEWS6bsLJEmqG
EDLb8RO4apKiv+BP1kMZPKamU4PCvGrRFnCrs93pCFiZw9ZjNXf+ryZ2jCbLYq3N2SKnRMrFQdYK
2Z6M9+tUypSBh1sCJIipkvkChlwSXVgGLPJtJ0gfPd1Ji74AYbG6nLFJq6QtePUuPqxbusLs9a1F
dxWmWlRfNX8N7j+jB05310GmysT5AYiNYnh/1oY2g8C9ZEkzEuBpHzgaxQ+Nj5JqawwRJtCEi6QT
ZvTXE5fMH0/Jb26SIQPL5dpesaZyjdJkpjO77ZUwouS3Ptnacawz6Fg04IJpjdkDjfZ2nk7i8n99
X8ERq2cx1qDeZbmetO43Fm2nBfkt7dqA+RoAccvo6LVmUp8ff3NmIN4i7hGQdkc5W39vjVAlNhYD
eXmPgJPhEI1F4Cxs5dinAfuAVQ4ZgiOD2en//+g4+zUSlmpu2rynTnwiB4nzTFo9YeyDIXeQeTv0
sYAi4xGWmxHvmpzTPvDRaXFU9Yh12UcJpWCMWyYG2pOvi1DY+ErFYCMoKASqLn3jIKB2XBQQxuU5
6NE7xXH7OKQ8L80HngE41Kdo0fvgTivQiKK8nPFOTErDqEUAe6j1JcUZEagiGPNW0zvS9LyBiyDb
jugFxqcq4d/2Vloh0r+l9nNSuL+yi+mJl9Rix0t2u/3+1HKtQ/7HMQAdlF3RwaVobHS5wzguYkUc
NBM8ODvbLUDwp7lmFaoZEPUkFjyPWDqvjuUbt3L/plaprgCUk4176Mv27EP5305OLGzDBYnHH/KC
CqVr+yrTX+yEGuLzIgi2CVw5RHQGXLnntSk8LmephgWAVQHDwGJRmOv0eUQWONDWFVteQ5eRmid9
9WNgeudunWMWlfATFpstJWt+mAiAcZZ5K3gUlmdj2fh3Cf+HJOdL78lZpQG6TBtxaR22xqUaQ5J1
DE7qcL7EGBKWMbIAziy0ZUcPZx1SC81OqwLtq0LVbviGSDTk9/MbGD7tFwlIwHMCTOqo4J5IsWQS
7MRF2RA7PJmrXM/g6Oq418a02Pat9a78V+sT+lSVrCMEr3zHJaipslwwgmr2ODodxg0W9S+ZMza6
UB2LnmWOzV5DTpoZpW8Dm73dYKLntr0B+U2pBvT8QbCdeU/HmNHfYXlCjQFIyhOWxrDohbEbrs/8
IraSgbBE2809d1qR3/mQwtb2hsMWG8Q5U9wdtZvA+uLaRCdRf0hhIBQMQP0vaU43M3eGygaRZWx7
bBki0Jfb52uei9rYeU0qvBe8ZeTXWEhhrIV06OGzrZD2QHfJAuBySbVe0joJ+YjDeyHvkdau/j58
tCPbKcEEhg9NSepyLZsZVBtlkSwAtyQ+AigKPboHLyGqoZLUN3D43MQYiOw6mMEorni4MQW3HyZJ
0cF4srC6jSFXqItvSy45fSbL5X0WnRNXCVHH1qO8bSs7zn9cAb8meIIJNrr1uRTELPXKMNMiVPRe
4jhLKCKvwpp2X5KxLHcNSC3lHTz93Jy5tY6tpNxUeQCRpYmzdpAE8jwOFZSy3Gs6K8eyS+4ZM/mi
+GsPkZ6I4KcvRGyDG5vTj0RQ+ILGiEstUfyo6Bex6qnXYYKghnlNgFbxDiAP/x2jj1UG9Tp1kGAI
fMGzwVbyBexyQ41iPkEeec5cictkhBdU0QI9au8fdWRZmWDsBxt2AW5/QeoXlxN1AxDS4Dn7yTUo
8BaPw+iDH7btgJuWg2A8jlBC+1GYC4Jj1vUFsoF+TuR6K2MIu8opm3u4tTs2eYBNIZBpAlOsyurx
2rTZMwp46ASwQyT2JnSNyvltuyCVIDbvltoexP7qgSTpXPGdFltM/BvKguVSufC85+iXFtP82VcX
+htUiTxyFuRGbcpwVO5q57b8ViLsRuvulwHloLguFk+gz/5Vfl84wWnIMPI8v2z6bJc3gfbJRq7N
6d+PfphwaWjv81i/YQBnXsLtKdlk2gSnrASGTn9ZjWnIdRgHjzfWvFY5wgqRRX2f/ESMLR3DXoDU
vZM1fpVqZqdKyoTxRCtU48eMp4UPLliYBbuVVJJR1kO+rmaLn3Yc6UbN71HKMilEddBpA6zFSDqB
kL21BYn7eAQ52CDOVrCisZsCP1fLQGtGzx/u6NFe81TVAzQcKktaV9NiQH0ZiLtlaAub7XcrJetD
1yviMV+i4dMuNNpLW2YGSgI1sNobosREOmsyn7Uif2zCNjJn3yqhvN8RBMFqstKM7mEpnaeVOn0C
1PvBEVa4+28F8KzkIRGzjgg7MAlHTuIvmG1s3u5ptqa2879WDla3cjM+gePPtxm1vafOp4C8fHgk
psqX3TcgQGhNiMYJTWxQinkiTSTcG6fZN+t1NG+GCheI7RP0q0OWK8H8M9OGmPldOR37zPQxpOjU
cFNFouDedOPHgdoUfC98rcuIOzRF5qs1mRozVi+K0q0LgZqazERWGqg9neT3klKQTG9EV17iNxZi
sj6UwuBTCBAPCsMEDB7h1ckNCnWIH/cMUEjQbTcFbvaZ8i2MG1zDxKA73l45kKc9w2uiI+nydPEP
BgmA32GbRWShTAqK/6s4JQpNWyrj5IjjMrXGG4hHDPGHRo0gw5WoXCNw/OBnsbaAgeV3kXsqhAYY
4Yn4PkF9eY6TtiVGDkOxgyfIPWVmpMQKmQUMRK4JEbg07hqEVvphe1utZXRSXRZV3RGxGxfk/6FC
RxPKL20po+J5mZt7zlUuIFORiydx8t2MjuvmpOGnMRpKIR0npZMjkwctJPX7eNZNAa+MLJ1uPLnI
fk4Jd4+I2XGIBTVuJrLL3Q05AGOnqpnVjSll9Sk4DnfauAEcQJ8Sak4+ZSkIZ5JLID7gL4IV2ln3
PFIz0G5cFv03AbBUQpO9bV9DsR9xGK7Q0EsjpGUcUVlMCaQWChB7I/Wd/YAqUqAurtwWp6YZi+hE
tzNqla8UV3q+R5b02TjhrOtzSdlGGNklSGfv+6fPsJDoAH2bXMmMWdB7LegKBk9221NvIzsX5t1u
PcRv3MEnRSuU7L+pgE5QF2beizR3PRaYov44Q7WLdhRWhQXrYcNAShx6+Juo5iWZmE2nk25f0GbP
epU8Oy1sTo1GPg0z6POmXlSRDQWthJYAYv9calfamVKPOgu12UO4W+4XxaxkHKX/5j3kBZKkz9YX
ChOlCBunY/MzvZlJ95WvND1FQKbcDO1yjy9AXvA+hLKcX0iuPS//afTjLTzKoewQAUZZXQoCJf5U
0rXvQVj7AIrTp9FlzPBUpyEzJuYyM95VrAt6L+p3DBcUYQ8QFOIbmtymyJGXgIXWkg+etYuVAL7s
PY/ZrarDOEJXtZdV1kQPCOrwAgiJj167SPzxfi6BJmNiazZ9dURpcfjNxPB7hNWJZezxVyoOOzI3
OGfCwjLU7+lie+rir5FVrpCOKVdyTaOeBb0cAcu+T3huu5r2kkEsxsgD+rd58ov+4KarvMPO/PRe
Yw9vdDd2+ZnbyUY6fOKDUutd29EjWxorMQwOr646E4EjOiiE3okpNR/PUvfuOeYLXWvKzHnw9gS4
Iaf1h8Vf9nQYCM8VI5hZiSu2t0slY14CmmPmyK4akQWr2MRbqEkVF6X5qFI24KjAW/jnQ/LX3dAk
0iaRtQX0m90FIn1/KMfoirhFkvjeHu4szCPZfsVVaNQB3xbSYoZ02Vxo94Q9ppnEVEt94bh25H/F
n3F4S5sPCruNStjRCtbdJQFMXH0nd3b9lg2VHLwK9Hh9hWCgwr0tjwSzuKiWJmcyEKXAhnE5fv8b
rUW2IkkPjbbJX3MadyTSFIOK+tecTU6hPXFm5eLOcAxWu5PrNKddzXGEjo7ZU4ZYTaebOv+bBtkV
73ZiHPyCEcVzxoAFSAVwBOkyQcsQrWLRZgBG3aCLVwuXRHO2o3B9YJvEywV3gnzcQi2ytvNP1cdh
HqcX5J3uu6wyLQ8jxtUZ0VLuSJUWE2/6tkzUe+rMo/yjiYV5NqjJfw+lJNT54zKHf+7oyHAbA4jD
o5YWZqei2LDT54bScprzwPuIgBE1E7WbLQNEhLHP8KIkBsW8dxM2OWIn26k033fsv1Wog6ElAIji
GPz2j6VKyMOMcfaTO0J1I8+CslsJppyFHKoxs5LtNHXrVAanGAiZm5xOx0SeEq9azsXF+lTPTCKF
eSDRqeVr2qKcLP8EehAjQpSrQ3oVcwdMEuiu3vsFnj8SOqHBeZWGvgQcfAdVgxMjTXnr6GCBvoNU
2gZoFmcNaJqCgAP5LoTf2s7o3R44lXSAnXvnkD3Gpem2eAiJAyUuNaHeDoS3l0F4d9TcV8LuFqaI
2JGpxWqq5KsjrUF+RGZXmyBv1hb9SulBjdHzcq52CEexq4wRAi+i/ugy/JKQ4vbrN3izOCv9fMWQ
ES6L5F/I80aKvVtk+1FdwhiK4eWFjOgOvW3p9Dalnd/eHj7/gJvH8ixL7+fcFqxkiZakmqQwP9aT
q+tDw8xBZb+izjs02oTxypn3An90BHt4/+NzBLTTGoLQA7xl7g4Y+nKH2c7qhImNlDryOozxFozw
yZVaeVCOAWi5BsJL35uo3NTKRtT7++hkvbLic0ghNGkdmJXHcXqVTdb5DH3oARH6IdyvTVEs1BLn
WsUTbRpbGgAv5r3N/H2rOe46fg1hfoYzCo+srDut3ZLMHT8UmaUlYGc8MpM3x7JH8WxrKK+C7iKV
VOoZwx3/D/f8Z8zI/qEgtRualIdRMJ3kkXXhmOZSyj+yTwS8vRPHOuGXVXB7uer2KhSUF8XifG8p
L8mgYhvsJWq4oeTxzOqcMpOTm6D9o4azAZ1r9+qz8C+FxhqLaCbv5KAMcJefBPiy3fxs78CB+qUW
Hs3P09yysGNOtJlFLEF3LHzeEg+9+kotAv78tRH+lIR8izDMTmNezormiswivo4Eh7eefHcyDjxf
WFVBM85Sz5aEe/75I8w15L/IhNhUQaOQVjTx0Gz5xEMnBarKoZyw9FBp8DfZTOsk2dm2YBJcuru+
BsewkhyylNCp6UBQPFD4ivBC8/8R82h9MvKqN57Rv5eDuGRP2zMMO5c8BqcuycyPBN2r9LF7gbCo
6CN5T5XqtSVxInV6UeAF2b1NL9qHZ2rw6UgRnTLgnng/Gm3cJhG4C5Z7S+gqPt9qcWVK4R3aDCCd
j9wb4GsoQsWVMwvUlK9qizH8ZhoZMWdgqnIsekB8/QsagoQlhsavAKN4c8ZXF6NO24n/pshueVlB
7Txr/gYRnZ3eiIqLqQPodcleqjQHpIT0dp1lIdZX7fL3lG/w37RAJxI3CtYOlBBxq+rHiJx9hByU
3HklI6l8/No/IRD+p1jAFFAKuETfba/QhNMvm+PvpSE4jn/Pna8u4b34D5b5PR+kD1Hk2/7jDz6h
Wu8IV/NVbp6jZ4b4vFL8aOK/pxvmLZjTxAE1UbmVZcyhD1xPTldvXWzHlbcuNIHUuTNeXfDqFr6H
g0DeWumzW1CmCoaWJgzrcc3AIJFWlGP0eZCyrGVc8i6uUM4aho+OqU+YO/b5BsF9Z83SiK8bwrRp
txYDU8U1NlV73ltjly2hcBddsCtvvciqQKct305ueI5pg/mdfiMo8PBYVi77NSCPCR8/rGzOMkzW
XecG9rcsAEG3f7yYXdT8fS09QcN3XdQ4D4+622FdQAtHgaw6NmE8r6S47zQzjYagSQ5N2iTbRoKK
9AP+trlbJy+gDAoxyUJ73NtomxmNLm1lkJjpb1jiImUogA2+qLg/cMXsJXYadhvFrKumGE8smd2Z
ztmAa8NVFOVDnNZ/z/BUSnjcnscRAV2g97dzS3czSV/5kHNoIqNjPxPHQ8CiZEJhCT3b88oS1aUW
Qju2EuBPhekH1Gnq6b//4lJENmstYID1ow4wHWoyYQQOflKjOHU2s4ZPa9FgL2Vely0TFC930dSr
/+TjMeRa3wwTy/8rH3FAUBnqd/uCIkHJ3agVRwR+T4lX5Mx3Nr6RxcQSLUjqFG3I4c2ufo5XMp68
hHt6zvbtyXT5VjWxubDQfEDUiJgByZemXqjWlPtPwux+s5r+/BBj1p8rKa9Up4NPp3coiVNU0KAG
zmQ=
`pragma protect end_protected
