��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a���V�h�x�����>�`���o��藶���ý�T��U�Sy���So�x����t��6T�0pnn,Y��FJ%
���t4��b@�3|�W�zR5M'�%�+�o\n��m[��v&��N���n3mŅ��}L���"�̞-��r��8tHY���� :�.Z�K���#G�*�5��s�e��gl0I��ddY��ܤ���?�R\(�n�O��6�*y$�����@����1Q�;ǀ�^2�a�Z���G��92΃ 1��+Zq�������N{!���*�)}�te�E��|�N]G*�۷t'M$�C_g����|�yAa�Y���eĥ���n���2�������(
�33�Ty�V�)+#���f%	͸4�Gp����v]% o�� %�/k��O`�����$��:/Mg��t����e�An�U[�D���n��X�|$�y~�͠�����e��V~?]g��%;98Sm88�NK���F��d��t��9���t�Y.^G���HC|��:�B���Շ�f ��Q��!>���O��Gp�n&�i(�ͽA��#mq_Cj��Nz>R_�R���׸q:]� ��VR�7�=ǰ�)�)4^�4%��>7��O���os�Y}������\#t���sS�2�"�
����J'���Hw�}3���:E���ޑ;�S��)�	�7�ʹ(�����}ƄQ�������������Pv%T���ב!�2�����6��`��!�>ӡ,�EΔ����D-)�o�ha+�"h!�f��uN��;����B�����L��_$�Db�Z��)��^�e�'�)u��/N���G_ ����V�J$%�x2��Z�� :�0��ᒂv���4M�Xm�+��[���8)!ckÌ#������`�K���B�5M�m`w�+��=�؟
+i���0(��O]^�;�aH]�ne<^������-|���'�ݣ���>0�FOHgk���
�[{�N�ˠ~�h0h�\ŉ��qz*Cu	o�Xw�pJ���9�W~�?Q�L0D@Q�4���,�Ҷn�:���Bw[�\�isǠlK���9.����6:��M��8mB��	����h�/��*NCG=�T�����ڌL�Uamt.������3Q�X���rkMQ�tӹ�`b����f?sRkcx�4~����x�@�)u����|?wy�uvX�˓-=U�`�*�e;GY�[�9uț�/�vi�(��I��hSFg�5���B�o�6%���R�@U�QeQ�D�q{(_IT��#[�7|l���t!㎍�y������L�N#�4�(��&���V��a�vp���{{����B�����6|��}{:OY(�;x�`�zXD,�x")���t32t$:�(i���׮��f���\>A �C�F/�+M���:}U^Ɍ�l!-;l����|h���W˜�84�5䡴-U��I�P:#$�ԏ�շ���h~"�Ftq����(Z�ՈZ�AwI���΋���jo���$��^�쎢���n�=�<L8�#>q}�����c�!���G��n��Z��z��E�jkS��J�e���J��W��x�$�	`4���$fX�s���
W~L����"��y���o���]�d�j�;*�H�1�zi�Y&����l<"[�|��<��Eno_e��$�_��4M����ύ���:�\�+�=�=3�~a�}=�ʸ\�\R��k�8�q��Y��C�o��B4��Drg�A9�_>�np�S�ƫu`������5Վ�N�me~nr_O������o1���]ok��t�A̕���j)��S���3�]m$F���ל#PXSi�ՙ�7]mY�i � �b�i��j*a� ���� �D�q��~�=x�E<H,��G����9 �ņ���9�~N7��@�}U����V��1����U��4���������l���)#�k�F�-A��@j�CV�-�����,�y�7�D��
��*W��Z-`���5I�h� �@�$���|͉	lkk�DE��2g�� �*wކ7�ټ�%rr��f�z��#�H�2V:'ne��}	ñ|�����F�$1i�!}��uO=�������!��8�ٌ�&m�_�v���ռ����!EG�3ݶ#V�Īю��w펷EY��U����o��U�����K��N��Ԛ�ڛv'�����\�E��ԗ�H%2�Ḏ� Uacφ�Q�����ߋPo t�)��<�>Ùu��n��H_��т뻀����I~�P�������(��T���ep.�rh#��t������c���m/3"�J�c�vN\�a��P�����Z��8y�<�E�f�n�v�tqȄ�)�*i�S�ԌGq %8~+�h�<FW[���7�w��d)����W�¯�x-��7�}����G���1��y�o�QS}L����6޸�"F��S��%[5�"��^�H�6�v��Rϧ������x�8~o>k�;��W	���ܣ�Kq��U3�D�#���_�o߾{mml�됫\�<�"�A��T�55�����kN�'��$�Vo.�]cG�@mB*�tWp�'�P����ƶ�2c�CH[�๏�g99%�Ǵ���sia32V�܌&����!�3�����J�����a!��A��M��R��*�|VmTM�y�$M��#q�.�)���R�-�1�����j$��HR�f��kr�³����	��'�]@i_w��o�7
^�k���6�$�eܡ݆k�f^Y�Lb�^���hyqFݰ ǰlT�4��m� �Eg�n%e
�7�[���!�]ā9B�m��@t�_���Z{\H�n<;ߝ��ac�DR�������h��ȥG;��r��4C��f$��]�,"I���6ecr+����u�/��_w#�t�����Ӟ�ԉ���ID���?���rc�H|�0B�,�,Ư�ۭ%G�0~#������I�dX�ޟ-Y�����o�K�h��E� ¸�K,���2
V��N�8[8F���q�z�)�DQ<��u�
~����]Ň���^}��-c�`H��Y^�������I�Kh���~�W��8eo䮽���BiYk^"	[r��m��s�t��#�:��{w��~(�0�Wh�?�]4���q/���ɝ&�� �@�zr"p�^0��0���_��êZ�w�m��c�i�x�c���(�,�X��_�eY8�"�S��:��Vs��C����}�����Ҽ<�^�}����ћ3�,[wH픉�
��@Ĭ�T$T槄��l��F�����TT�2��q |��:^�,�F�G `j��Mvuo����n�tN�L��vۂ��Z�PQͬm��7�l�D�=�[&��.^�v-����P�؅~[�LGڃ"0���.ag�C��6]�������R�����F�8�s�[�B?ݘ�����"��
߿
0���e!h�fG$���Ç�ლQ�9#Dq� �������P���s���O+�\�6߲v'����r�&������P�OuoVU*.ӨBb��ެA�a�� �d[�+�k��揭�z�6�y�K◎NW����ck)�TR)��av(�o��-�}8ć+���%�L|����9Z�O\&���������]�ʦbNf�'�k��cJ
D�B2��ڐ+�|�r����N�r"����f�k;h��
����8�����v�I��c �D*-�G����v�� o��z�\,7L�$��r���|N),�N�7�b�&?0x��A0��#�i�.�R�����ճ���������KYŒq��TM#:�o��J5+�6�)R�]3Rm�I�>����"��#�II�+x�F�ݚ�B��㵘m<��fQ6�^�76�>�`P�C>j<�noΒ�,���h.輢�
kGY�ʍU��/t�(�c/X4����B����I��}�[iXl�jA��?]&���P���P[�?�/"�~��bBrT�߯�a��X�Ɨr�za��E��Ɍ����E��b��XB�o�B�	�`<]��ŵ��KH�ZϬ�=��������-�\�.;;9�� ���h��8�Ks�H���6'ڜ�w�?g�'J�v������,cլ�X�%JN��nlY��c�c�)��)ۣs�5
����<\��G1���0�kI]j6��f9O�Զm�}�t�I�ƀ��4S�	ࡉs7~�#ɬ;}��S�}M㘘�C�R��Jg��̇�� ��&Z�fwy��-}!HU�E�����f�YuqfN�Y�����-��5݆$h>��;	ZL��1����RzD���� V�L1)�A٬�-6Ro@w�����`A�T�\��\�L/	�yy���� /'0�FY�r��v��*#s,xy�����y{ZE̺����a1��W��b�B� ��1b��f��jp��x��T���*�_�&6l"q	G��-�B�.?�&TLP�ٝ������M��Y�t��tJ=��-�f������Z���:}��?���ʆq���L��"�
`gկ��h4�OxN���q�~Ο'H��~Yt��=��\`"��{9<���FL��-���Oɞ�Q�L�J�^u7ҵ�#j�8��j	���7RK� q�k����7̍��%@~�w$���$M�ߠ�s��w�t�M�����h)%��Y�)�t�W�l.�?�pJ�>EZ|���jG�i���[�wƕM?E�b����F��`�y��ӡL�ޣq�%<�J=��@A����:��_���@X�C���0;J�(p�x�C%�fY�N��'}��T%�,������%թW��yƾ@{8u��<�7[��d^�m$�*�����0��K�0�tʬ�1BC�:v�_-�Ӕv2��p>������c�����'��Z��X"�_�}��I6��\�^P�"�s�DFCv��v��w1s�ߡ@���gm1'q�y�!/K�=�E�y�!�g	��D��
w&zVu=���:�ԅ#���o�OEs�?U�㜶��;�r��L���3LT�D��6���f��-T�.��з�F�<��GyP�į�T��KZt{Nnc�NL~L�f��y�J˽���{�~E0~�72Hd
�,�u�-{�y�W��^1M����7._��Ԃ8Mk�xkB73@<��N��5���r��+7��+��N���~�D<�A��qd�>0Q~�yZ��f�` �-ӎ�m.�P��+�4��ᬄ�����r�ho�f��ˍ~��#Q�8fLº�dW��w�0I��z�Q�Â ��d���eD��c�����歧r�����?��(��ˏ�}Xi�q�H��$�ᦗ�?;�S�%�*oP���C.w���7��j"V�0��N���*�u����eA�7X]u�/ܬ)֬o�Q�` �?��9�t�{-L�{���T}U�15�ۯ�4�����a%�k[�2k�G��Ʊ�l�A:B�[FC|����c�*�-��M"�x���Y�����6`��l�3�Ђ�I�!D[��͵4�(bt�R��.�D^H�ۤ+=��"��D:�輩{=�6��N���,l?o|�Oco�l�i�u��"�^�Y>iE�� �uV�[U)�� ���n3�)K�":Eę�C���WEa��HN~��Q쐓�֝1��#oZ���$s(��Ҷ�'�%�G�E�9��Ѽ�b��d�ʴjS
C}���3@�g��:rf���ɰrǀc���R^w�u�I�F����o���#.ӠEj\.�ת��2빮Qr������S�;��
M@`q�~�Z�f�Y��������E� ��8����Й�<S��xw�ۀ0���W��}�Y��?��cnSQ�|)O��]��$g/�3��ۣ!=�0�2dc�A�f��l0�Z�\3:�.!ᣕ��\��V���Ꙣ��2&KGĚ�(ߗ�p	��Ɵ!��:Da��8�¨Dg�l�g|V�4�p�lՈ�(iQվ.�ч�(�ߝ��\�\�]t����%Ƌ7�g���DAE�+
aU�1��꧳�8'j�x��T8v�I���I-;f;���e���cf\G��J� �|_�,�%e7A���adgٍ�vx �0��)o�Xq�m�9/��{�}k�1�{�.�5�[[����xW�$�6�~kC���ڌ�Q�	?�u��'{�Ɩ�E;�G��>"ɮ�����,G��@�/+������
��$��l���ޙ�Wn�A�_�X�3�`��K�:VO~ɻ�+�� 8�Z��y��Ｆ�y����vcjSa���'Eu�A��q�@�1��� K���yC+/"�e�Eъ��N!�L�2��g�Qy`�Z:�����ٛ��$q����arh�"����V#�@�[6��µ:!`���̭ɴQ!6<�����	��i���<�!Z.ӗ��N�k1?��q�_֦�c�v��l�`��(Ȋe6fj9j^����ƅ��5Zf�)=W&z��f���nPgttZ�=�����r>�cl��z��׳��e���3��ԣ���_a�	Qb�5jtc�A���G1
)2̮� ����+�Ė$�\�$��:��,!Ic������s`6�c���dC_����� /��3{��V�Q�f��Sw�޼�{X�5��b��[������}n�!B���O��0=���Җ]f�K[H������_AA��j[��4xW�l#,U�R�Fh��Z��e%�Z_s�A��V�I�]�#b̖��w:�tYy��ոj8Z�Xu�J�?�S���J��H�������8�`ޱD������v�BJRer�f�e�O�;Z�v`�*���AWP3?���;0�:�����U4HI�N�1��r��0_���I\�E+X'�w�X	&x���DdF�X�5��< x�d4�\�H�H��aD��v�FuH6f9�:�j�܆L*��d!����F��Ӹ]��N/�`�P5�c ���k���b!���������R�"��,�ϋ��R��CX<R|����*
�S��k}V&�<ν]�+�֗Ãme�H���&�5fy���hdP>Jɹ�$F�dt;C����5��� �F
%vBf׃
]�;(�`��Ihi�%ǹ,Jb��?3���d�g���;�~�o?�D���x�����k����c7����\�W��١&%��<�PJ�ҹh��b�I�[ꎗ��'b�����n�Z,�[�\~�~]^~�#Ee��5�<zH� K��Nx�f�&!t��s_n��0ۀ�F�)�/s5!�B@�����F ��U��qŠ�k����r���±�#h��!rw7�I.���SI�?������_|}������u��#�:0�_� ��]^C��͖~�&e�Xbv-.���fm` ��qkؓ9S*�ͧ�ef�0xu<|O��" ��g]�s�p��T�WW侩4Q�Co_�毵;ǭA 3��=}IC\-[��rm@���:�Xa#�%�p#~.
�w<��r	���� ����y���TF	�����a�^-bt����|�\��H5��խ"$�rx!A�P��z�Z�1��H�ԍ=z$��A�"O�f�����n�:�Б�܊��`b���m �����;]��nb����l�%���;_d��ޢ��W��a�+qj�	t$�[X�Sgd\�'	2sB�{�|fds�����A2\)��R�M�i�y8;P�f��p�a�Z�S�wt&���
1+'���ⳟ��_D� ���ҏn�}�C���b������$���m-o�ӛ���'�|Z_]� ��)�.����׷ˀ��>E2,��>iU=�1�tט3��x�+����cF@��i���������-�G^,�<n�,"AX�#�1*�s�������D��Wꌒɳ���'n�� ���`��R��A$�s̑ �{ �_�<(��2�yɂ z�1�;�0��{8���L���/�;���I�Zl��C򄂟�M��> �9�S|�I��l�!ej�q-��y��� �R�L�/��؊�Q�"3�@�y���f�b���3�1�����2s�Ӝ9�S��?j����j�jĞ�e����KC�e� ]N�z�L�*I�J6�
��h���]�B����q�]Vk� ~n��C�����|�zܽ�C&%�+Y���µ���ln_�G�S�͖�֥��+�V5���f����f�p<-��~��1�(��W حC޽`Ori=��a�`�O�Yyt�Z��^���пD�:�͗����Z������ΆLU<������d}T�\���}f�"�ֳ*g�sf��^�LŸL3K?X�%;0�x�,�K��PyU�]�\�|��+�z����d7��Td�9��5~:�����Ŧu=s�r����t����1�	H�ML�`nm����&o�c�<U����o[�V7�x=:t[)�5��%k����~�u�����Rf���P^���O�3Y i��	��ҙ�����,Q�.24A�.�}��)������]�9�	��ġ�,*�e����p����(�9b,F�{��'��<|Pl3�s@�?RiÚ�n�L031K�G-1�E?Q�z	4�,�`�>�I����6��Oc�ԯX��{Fy��� M>��U�D�ҪZ����K߬k�d�acy����l�d��b�B��O�\���K���Eѷ��_G4���2��{~�hE�d#��U0E`'���_�u���Y��V`H�֩� B�l+���de��i�����\�Z��~RvO���>�,8k|ߞ��X�y~��i�!��@��3w�]��C}P�٩�@
#�����r˫ŗ����W���&PW���3:�_כI7{8��io5%<�}�P�N�<EA��=.N�<T�q'�V1�[O&	�ƴ�B�t����]�kF`��-&�9<�A8|��� $���t$~�H�.<�G���`�'�B�G�_P{[�4�F�n��t�b �Z���s'������(^�P$�]�@�Y}{�66��#��bȸ�ʶ-��[�Kp鏤� 04]�g�Vq��BD��pC:+N�����i��YG ��̈́��t���%Ʉ���q<2Eϛ�S�v��+���<�l�(��K����k�!�9��l�a�"+uM|�ٕD9��.�c,��h�y�/�`psu�v2�I⋔8�3 �����*^�G����� �P�3Ă[`�J�&�Lxu�~W]}i�А�h�+���� n�S��~���$��XJH4�ǎ��g��v��w5p�N4-�Y}�"S	�5�ZL�X����fУ:�	t�0J$L�\��9:��i��oΥ��0∛T��ܥ@�mp�aO��aP�[ ���.̃�.�7�|%�����aBpE��FP)�y��YøJ�=�h���6��we��D2^5��������xg��8��؞�+bG�U^K�w;)Ig�!�D#m>�Ɔ���1K����=+�'i�`|�ך
j/����V����Q)K�JXUl������~36���ߴ�.���1��LFp�����$0�]�\����u�"�R��j�,!�տ�/ y�<�p��@��oP���.�8�;�V%&�u��lauF���y��w�VI��4(
���gr�7��2��y$`6�Qi��x9r�!�]�CG�v>N\S�P`�(�Po�����ӗ����������}�Ɲǟf4v�n�()�O�\-��v��mM��I�	qK�4dX
�"��Z�ěDDj�J�Uώ�����K��cd�K��\\`��Z�n� �����5����ُ��?Z�N��'�7��i��_s(��*��WCq"�g�	���-����MI�m\f+VC��x�- �&��>���,��9D��)��o{�����T�=9�Լ��F�Ȳ3�J��3309��s'��dVEY0s�yHd� �2iUN��>e6*-�(X�:��w�w�>��%&��gP_p2Q3e����B7�3۴�_7V���d,p��Sj�4= 7j��i���=�7m��{[
�Ct�[����̇L��a�-��T�rL�T�s�ú�X�� �5g}.S�6�.�O��C�����e�HOwO�>��5p��������7(�jb�5�v����`�i�YJ��')�]�GkZ�u͖b��<���5ϑ۰�.A�B�G�����$���X�`̹� )l,�BU
H�y�����S�ڏ>|�3�2Q�7�Ӟ_��{��(Ghp������}� t��A���o_ b^����-��8\>�]
sI!�
<M־�e9põ1�|�fؒ�a�oa:������͔���G��ݲ�R�c �B�y�����z�y��u�>�0;���|s�R��a��A�W��}	�;։�vU��P`��NwU�'��}��W�������]�-B/N�,�yF"�|=�S�8I��H�aCt��-��KqL�'RB�������i�����n̗7�
H��S�;�M���%�2ߞ�ӥ���5�W1��^���?F$���b7�P�'���zrA�o�m�ށ���&:�@�k\�%T��=�%��B:�����Olz)1�� ��̖!�8uᴘ[����Ĝ��dٳT$���.�k"C����7�~�h�N�40|�%������>�R�`���@��RME�C�"�Z�S����hF�����X����+�x&�F�/;�Y��7�ޯ��	<_^=��-Fe�8n�Փ�jDL��_��md�#6���o�r6LcO��?Jp�>+���8�:�pI�K��#���i�M5�K�ip�|!M�4�l4�4�ا�xM~�GJ��E���wt��6��	�/�@n���^J(	5��nd�lu��nK}�4��y-�*(�2J��|����Ǣׅ���d_��A�#�΢EF��~3\�*��{;�:6�4�o����gD�҇����O��Q���>1UG���78�\�+ьh�?`Bc�m��φ�����ŬHc��SǺ��@�����(�8���G�u-A�!}*�%����Bd�V��%�)�s3�u/�d���C�%!f���肠]��̲�~n���܃��e1��		����� 7?��PZ|V�����!멏�V���`҅����g@'�}ύ�4�My���	�h&J"�YA��pː�:л"4� *�]]9�4�+���\���J�I�JMȅ5Z��s]��&�e=��o����2Z�pH�"���ߢ c��ٿ�Ow�6gEٱ�l�Jm95�Xp���d�\�cC}ϭ�iFj�+�����Ji��-�_	Z�)�ާ��hj��dU��b4��<�{4�6�B����C��hs����x�)]ߜB.)L�$a����	�����צ��\Y"w>Ɖ�\6�	���\I�hO��:J?<�1ݾ�v@���VNc��ဿ�O�2VEa��	�H�[f��<�낓���M�hH5(����.�����5vR�I�9�rb]��2��'�j�X����P̓F���3L�׊hO�.�6����ݹ��Q?�g���-e<?���F��������$�7�#��0�1�SV:�*��ߺ!���PP�Iw�!mŽ���3�q,�g�Tے�U��|����9L|څ��]G����q�9nV-�$��RB�4(k_'cWO���(�g���S(O�>K�=�ĸx����zi;�tr~'�F1`7�!��\�����abY��ʙh��c��c޳^���<����#���";{-P�����>�����_?	�i�k������h9ᗓ�s�Q�7kԏru����1�Vt5��ϲ����:�>��K��ܝ�Iab'��Iq�"�O,r�2��4�s����,{y���]X�xo��l���R���o����|T��7�]�p�g%�*I+H�����%W?8}޾���ǋ�Ύ��Tv���Te)f���eץ��j/��^�y�?U�){v>�E"ʯ��Ge�D_=���>Q����eo,f9�;�H\
��9�_Xͭ	S��I`�*=�
㞃mJ����h�na�y�aF�~*i0��IF�g|T�y!K�r�0��SĐ\I	����mnR|��E��b�0��'Zsug?���ε&ĭ[��_�����txgn��Y��}߳?Hw�ɦ��|W��t��D��N����c�qY!��t����a�p&r�G"mKy�~��攅H�Q�Bigٸ�Jߙ��N�7��R`�(�K�y��`�뵝�l��!�|��MH"?6�{>�c�	����� �ʉ+cX3�z}��ntc{����%l�j�t�~zh�\Ѻ�Jq���N���_�f��{��>��P�IJ���w�T{�:�o�/�t �-pM�������^&���>�w���/�*�l�m2��'���34* j�M��R�@6v���e�������6q���3�[x2�.���s�|ߠ�.B�[eK��&�8=0]N�-�����E�0�B�<��!���\�>�ͱ�Z2�ن��r�@�7w
2#F��`X�Uc��X�Y�����A���b� �$�,c9��:����P�w[�6�:q;=�\�hh� E�bɂ�<����ѢC�%�D�>��G9�U�ʆ�>F�� ����MCi�`ۼQη�&�(���q���?4�H@�H�.k�� �/#XYn�-(�@�
q}�%zQ�f�W�^XDe��_��wT%]Lfg�"!��th�ɤ�:��ZC�������{�o	�\t
D^)\��r3t��``4��Ad^��L��d_u�ʾ�Z-dc�h#C�pS��ԏVD(m�65���yC��锊ˎ~�%�E��3^c��ߐ��?,�˿�bغ��C��TaN���~3���oR��1܊BC�)�a��ܔ���^d�	��.����J�]Ң�N ͱx�&}����I�l�6��X���֛�%���GM�l�0�?��.��d���BA�,lJ��[�`G	$[�Y�7Y�$�~�kt�K"����R¦�e���Ã���]{Z�h���N�3������<��k)�����ƯJi��	�),V��p�r��9��򉡆��nM�[��*����,���A�[&�~�6/c�Fѹ}4��V�7
6m�86�t-x%4)t�P�3Ui_Q�9��yV���{�[/���hl�uJ�%��ѧO;��M�|�a�99��V<�K�a�t�����8�cb�d��GSZF7��#%%EA���R�ka�L�4T.��¸5[^R��ͯ�yx�	���ϕ�}���!�#��JL�K�q��QMc(wj���d�6!�d'��@MgBgD9m�E��8�z u�\#.7��{�=הT�MR���;�p@��߂XX)�Q����}��#-b�u�3���#YQE��acoks��s���{)��h�<��>j�Y|����5���E��*oZ���E�:]]�t4M�bn������ ]j���u�R���_?8b�U��aSB�OlN�զ�\������~�*�~K0�}�a�)YU�]���B��%��x�B��U���������W�UP��|�!��>���Bo �F�ǃ+��;�ۤ��uRf#
4mvUA�ّR�?�"[C�>��в^
W^�n?3TZoR�iS	�>����T��F<�c�6KUK%iPM[fdv�"+?��qfI���q�nRXzd����4�Ä�T�,���	X�%�RW?��G�)N�l�W��DŰ������%��X�������㡆{vw�Q�!..�%���D�p�,9i����'��s��h<d�������ɥ{V$Y�{�h6�K�Y�$\PAt��\U�m ��4nd��	gud@e�<��uA��'�e�+T�M�U���L$�����5*��!-�6rd��юkֹ4�P�� ěY��l�Fb��,��,�˓���`tdJ���Ҫ���҃����q�D���l,-��Ʈ�عU����UVo�D�����ew�J���l��)
�X0�S�Vp�z�6C�����rq�Gt�5L3<͉m�d�i��ᴋ�y�,>L?a��O����-&>[�)��t�Q���+�}�������!�;3�����y|��4o���!�,�����&��b��OsX.�G;�?���$3�96e5/9�lKO��-C=� �q%U�h����	s-�8x��-"�k�$��f������G�78�q�=J�)�q���@�^΁s��շH���*}�����a��� �k���'w3(�2�%��v.A0�)��O��g�g'��Q���X��b��.���=Ă� k;��B���K�޷���]\���z�q�������n�o~��V��o�T�w Gg�Q�u����@,�#{D���mW��6�b9����u�����r�j4�v�8�6�����zVm�A�>
���#�xOj�� mZ��(���lUuy��us,aj��K��x���2���������7��j��m�}��Z�D��K=r�|8���#�.��a-pɘlՂe ���ж��:����\���C�|%���	���5:0�]��	�P���np����}ZD�	R0�DXE�I��<-f�M���c�wy0$������&!�u��8��G�� ���#\��?MhP����u"��r!�a�.�	5�u
��,X� R<�ɸ���>#F�N�&M3jk�����#2x�K�@z}8]��x ��b�#��I�UhCk��+F����2l�E�j�3��[m���-Hoh��5�%\ԏߑK�e��
^�qaEB�-n�M;��r}��)�dL���?f��������xdS<'d.]�]��E�����bƧ��`&DW:�]�����`��G��%�(���*!xz����x�P{����o#ӝ�V��~���83���ɳ��;���hm��=(��=\D�pt|JzǾ�D�v�_������Y�Q{f2|�ы�w���jt�UJ�����s�����FZ���/dFϳa�����1��7�^�|����I�L���ދ���m���ďmI.���cQ+U��"\M�`���Y��p�"����"��X*m���Ӿ� �	�����/�s��w��-0i3Y�Wh�o���(Ao� ����]x����Kr�_9�WCkW�8{��2��.sU���}yl��ݴ�Q�-�'�f�b׃휪X��߿:�����4s����y�S�UI��ઔ�f�u8�;�ļ$��~hai�9Қ�+D��~�V1Eh<e@п�w�Må���s��G(u�� ���U������Fo\��*ŝ�e[�4�/2�1��_�Soϣ�1�C�q��o��ˉ�w����X`�_ô*K�16�#�'1����ª�Fv�ڒ{�!I;U�O�}Us�9k�����H�T�H��T.O���A��i�J�DԽ%;��k8ܾ��ʗ5��o4E~�-��}g@�� ����'���j��=��1�Hi;�EP^���o|e���,.��}��OY,�FM�?z8�˶�	�|����;7I'�#2�4���i�+��]�il�N������)s�{����qV�͸F)��B�8�6?R��
�F�Jg��H�(s�r��+�KM��"���vH�[��V&��e��,���.���0UA L���o��g��$&�g�s� ZXcڅ�鐒�vP�ֿ�o�t��@hDLs<V_���8�m#1�����W7��0�4PmE�E��5{l���s�M3c�S�%�a�0�����q!g(G`�C,b�#��.�����W��#M$J�U�R�u�|*�2�/�nb�Τ�o�
����@#�:�1�8�M�hV�!1��m�/���p�����K6`��v����8;jh�b"�U�7��~��G��V�V���6~ E����Y+wÏ�ڂw�J��u+E�}�i"I�$zd����}�����P�J,MTK���=g:J&���Cȫ���,d�)����}@���J���-0�Ǉ�f����*�W	����RD��
���F�]n��t��ď�β�)�쀞�j����9x.������N~���~�P:jo��OP+n:���M�$���0�B�T��*!�>�rP��P�6J6�P8���%"��[?R�d�e��&h8�ip���J[l�N���K�L�
�4{����/�����E�^z߉�
�%��R�P��j/$�{���f%U�n�nf�������dGYm�i۳	�_P��.�R)#��:O�	�_���J��mt�q���j�a,�R�py ��d���E6���p�A�Foa��~N����*�׶��8�n1d�u��m��sy�yM�u�9��8r'�w�-ς�2�[��U�!U�"�#�l���?͋�sj>�C���M�F,wKΣ&!{���y����N��q�-����+�#IOk������+����Nƥ���@<����0o��<Gh�3Li�]����Ć�u\PΩ��{~�eMs`%��=�&v*3��Ue���w�Q��n�Yt-������#��T�N���(��Q�/�\���t�����}�H��\����Gq �$��Қa���R��o���'M�;�_Ԭ��v.o�����7��$�/��oK��=��l���ർ)$+�5�c]Ђ˅+�?���G�S� �bPf%�����JUf����T&�R�Nϡ���b�v�˹����3�\ʙZ�w�-�e�����P�S�r�{�q?<��\b
q�a<�����s�{
��X-q�ij<B4�/q
���z7��R�����4]���eт�z�����}dڴ�6/�8�-A/��I�#6'gy	"h�����]�)dm�pD�B�3�~���L̴�"7]�B�2ǥmW�X�t~�Ypao����/|}y k崗��3���>Qּ�yi��}��ʜ2l���:���y#���f�>�}pL���Ѩ��>�A���`�ɝ��7�(|��t {��_��Ұ�2�Rĺ��0E���s�K�	����kmq��$�á�����a��]П�$�Ќ�l���4�m��K��ߞ�B#�ԛɞ����W����{\�Vә�S�r^x��S��$��zt�@��J����ʉ�^�I����B���M�� R��#	[#��x�dNٲ�y;�I�G�A���8:x�u�vW;��s1�ĸf �(��c5].�F�M�?���)j���;��]�)�1�3���������`�Ղ��t���������ߗ��SN_���kP����]=��Q�����A]��Q�+�rz������1��|��ؕ"�R�,W/b./��=*zPr:B�Ǖ��R�,O���7�T���w
�'nPt�5!�蟅�S{5�@��=|�Ĭ6�������b��}�'��Xa��P�i��d�Xjqz�Q^�C�"�:�n2��X���X�n
������
�q{7�A�o^��=�qo'�]�T�w�yK[��be+5S�%�9Қ���~d�����Vf&) �AY+�I_2��S�����5X��^T�綉�+��ݽ��²b��!;ʒ�.���	�(����$�s�A�U!�
#�6;��"�б�c���X��fa���v�������\���{�ꩶKb���f�VA��AJw.Ls؄�a�-��gۛ|�#ܟۀ���&��ɵA3��9�,�D�R����!����j�Wl\�Q\������X��F�! y&!/*s}���jVNwm;C�
rу��ѕA���O����x;B6�a���c2\.*�=ǒ'�o������S���I�D8�ZN\�7�$�6#��Y)�*1u!�f�|��H��&o���9���?7x����q����$�̆&�,q�����5, �^���@?���0'f�bS.A�i.kg���&^�B�$���ʠqX�_�{`�-��"�M0$��Ve����AղݦRnԢj�$"+.����c�
M���#� �w'&"6P�Li{�p8��y{E�C8K������+�T�6�p�`��JE�4"ü���S΂|g�y$���$'	uxʷۑ�]#׋�C3{�
��DЬ���D����#k|��o5���'Kd.�R�&Ac(-|s���P�;�|?�ם\��Bwp�~�����IJ���Q�Ws��ݽ���:�>�ߝ!1^x�RH?
E� 2w*�ʢ�O)n�n��>_�-
��Hb����=Gb<0E��E�M��R��R�lR����#�Ю
Ŭg�$b�2d�jP�:VM����޺b=�'|�)"ao2�x�:h�V\���D��qc�����D�bc�����wp�E�aR���hT���x�z{��x|s�aW���|y��ۊǆ�J� �F	X��P.�A�,��5*��t�6�i�p�5����6�5�1��c/ͻ�����$��^Q�.K2���\�̟�Ex��e���{�,��]�q��VX��5
�����7����*G%����Fk�-�y���	�Q�?���$�Q����h<f��A��_N ����O(0��pZd�3M2����+�I��6��^ �9�i2]�����B���E0иB�I��5ޛ*� ���;Fm�³��"�!��w<���46zot���6?�
��ޜ�>�1yF	u ����>+�#���ZE��#aㆱ�����#��YB��!gG"1�Y#���X�c\�H���>�sy9�dH��E,h����ty61��8\·�y��c�X3���8�t�1�|�~M˚x�0U�ݴ(�s�������/?Uq�8�J�T�5u�GW�C��ğ�Jf�(`�D��]�md�.c%&�(�a!Y���VL��`�J�a�H�
T8���k�0c���_|K����]��p�&BG����	��Ҵʄے
^Rv������Yr'�y�=�`=L�vy�~����P<�)ۆc/�n�gv�n�|�1���F�"�lf�K
ilo7��aKj�TfO�D�|U�j�ȗ�;�Q7��2h �Y:�ƴy��9Ȟ�n4����N"���� �8oN�e1��+V-8�Λ���|���vZM�	*�MD%�!��K2p�������rzߒc���Ր�������'�ж\�Ə݀䟛�e�E0]������HÌ�BQ�2��dz�����t҂i��x3P-�z����|uj#�Y���`����+&�}l=4��Lղ��_�Ov�C���v]�W��_�qsNjt�4ԐuC'�+B ��R|�������aCEW<�}U��  �Ny�F�w�[f��L|<[�n�-	��U�9vFxH����u�ʍ*B��Wϡ=�ɪ�c���o��^��.�4�V�������b�yT��難j[���7�d2zS:
�6(��[��2uxQI�n�m�kR��T���%X���N��&ax�`�&��W�&�ŵ74�h��f"a�Y�Ho�؛����vGsK��b�\$�b�<������{�����YQǙL�~�\�=	�٢�����}����)�6�JV���Y^��x�Sꥣ�R�;���]l�<��=��]T�3��Fx+���Oח<��d���P�ۘT��m���~�W��5����Q��寎�ZŖ���7��c=�;�x嵄������~����W�8]ux�0�Ύ~��K�^~DJ;#��RQ�S�M=��I3K�����F��B�{����k����%��B�Н>��	
���;
�˥�F"Hҫ�Nj�����J��!K5<j��J�H�L�HŬ�R��@�O����+�v�=4��N0�2A�����`,�����������QQ��"
���"&aM���Խn��/��Kn��샔o�����Fr�5��-���p�x�Ϫ�Iz��%�7ƭ�۲��7��`E����6�'�P.,�xgB�`��})�ۣ��d�hU}�ߠ�	�A3h�g�J�̗e�Y�T�<r��mCL&�������5��kI,��]	#k����_�ēM"@Z��A�y�_R�)@���Y�Dy�͎�a�"Wߙ:��s��X�$CЮt�9
R"��G��\4۷ ���H���$jL������sh*@/y˥P���xx�~�O�q�� V�A�8�#�U�.�%�^���4�+���<�6�g��=l��]�H�Ճl�G8t"�[_m�+�Z�kNwh�[���|��u��q-E)���4a5��m��b
�g��d(�Z.��G<�-��Ũ��t_��.C��Ѕ0[�-����}$,�F�]�6�M�rm�o��T$����l����
lQS���ي�bF�R%<��\p�-�8%��L���E�`%%�g�n`�b##��x9���j�#=u$O�Z����[��?JsҀږ�4�F�.2j0j����ɨ�ozN�Y�ox.C��O�x��^Y�׈m�o��ևK3����|t�߇px
�Xbl:�������� ����Հ,d )�8����(ح����z<��qs2��W��L?�W�]Q5��85��'X���$}x�?9fߠ�3��q!^cf�EC����l�]г��H���'A�WvU�͖��蠠:�)I�4�gYC�텕�ο�̥L� W� Ě>%슞�[��s_+[����$� q�AQj�9�%����_x�x�}IW��c+I�i���9��G9�i�h	5�F�ٵVl�v ���0�pF`����To�f���~���K�ƭ'c����sV�iZ��*���9J�Aɢe�M��2$6����X�<^�'�
�}�H���=��H��_1I=!~�'Wݒ��&�\���ae�����h�ܫL�F�\�����ΜD��9� ?�`\��lyGQ��r{-E�F�q����0T�9��v�7�8f�	b\��sG��9dH����,A.��]�-y�Te�WP�S�ZJ�#Z�^Ox�@e��+DY�N~w�V�D�L-�<�7��<���L�UUU#Jx؜ۿK̬�����%ޕK�a$;*
�yr/���f�?�� T�<Sg�"��['/��X�ս�Ȼ��pdn��/���ג�#�З�6.A����#>�C*��ѽ���~HM\��x��e'S!��������z��i�ô��9�]����x�����TW�y��!<�
B������؏�5]�/��Q�b́%�)X�(��7=V4�!��T��4��ieDE=��M9Ҡ�����8���y5���-A�\�����G>�_|v�P��>-���=��G���t��)��Y���Ѝz	��� �^_{F�Z��1��������j���<�k�d�})��̅�#L��m�,�<��8��Â9�%s������6�GdIɐ�������L� zZ�Df�Y +-.���%�2��N��$���W�w�~\�����4v��Kw�@ۚI�!Uz�����*�eH�[���`���&suA��!���~_�ͬogi�+���6����~}o��J�w���܌��H�g��ŝzY�d
6�kgY�q{/��[Ӕ��I�����g�q�p�Xy!{��aY*AtW7[E]��@)p�w��U�ǧ����P���;ئGS��~t�"�"��t�d�W��B�̄uբ~����3=�#�ee��4/�{�"�*u9�B�ɚ�MHT�|Y��ɂxt4��ȋ#��2($��� ���0�ȅ� ��~�K����;j��y�,!������O��J5Ln�ʝq���	��Y�UyWm<xX���܃��>�>��m=S8�m�g�=Q�2�n����eX[v�DL�DʀQɊ�12G{�XY-��qS�E���%Đ�22Tp�My `�s�q~���Қ e�a�᎛m��݅�h�:��Ź>\3H`���z���J��~��B"�)Ծ���
�[�>磉�e�t��hZ������B�l9��NΒEX��pO�!���R?�!���_+P�l�b}����}�NL�p�	��z"��/�1����'�0��QI� 	��Q�:�p<���������B��5���IűJ��J�+�������A]<=�C8�>3[<�ǫg^�+�v5u_D1�F����zy-�}��#�>˽b�X���&��x�W4�s%�ְ��Y�����U+a���n��nq#E(ˇ,��e�F��Dwby��E���"��&|�?lpܿ%΋��WxV�/&��8�؛[#Ip~-r:m����b�J���x��>����e��Iz@W~�!1��ET�ܹ�v���]F3�ߝ��'�]�D�(�ͣ�r����$�G0O�Nn'�&5���8�X�I�Z��opU��z�;qNT�S�.�#S_D�g�H�l�^��7�Y��;�"b&��0����s��y#c�`��s�,	�-�����}-�����;|kзC�?V�B}״��r���:ƘF�`p�:d�wR~
�u�/�ݍ��9Q�+�|_�ڲ�Q�������l�~��W]6�jJ�(Ud��׍޶ٸH��B��"	�=�p�ˊE�5����QD\T�U*t�����A� �I(��x��h�
�+����������ů�~j&A����Ae�l�P��K��;Ҕ7����pz���Lu�׎�3��q�:P�:9毊�z/�A!�J����33P=ػ����Ւ�t�I�T	ݮ�Rx�:H���˯��G���@���}+Z(��u~ÏI�:��#�FÂ�U��ҹ����:�
a[&�ē.�#��&	�[���nl�����D��eɆ�QL�c���3�'A��¥���m}�$^��H�*`�]� h~��C�,�a�z~�Y�,:7��b/��Y�ʇi��*QX惟�;��(_+����͠a�q�刻/}����x������ս`g�(�.� 77�=d3م�u
��z��^``"lÊ�h����d-�%|Mr��4�K�@x���t][+{� ].$�TcP,V��>��Ė-���UP,��?��X;L�Ӈ6����r�Z��h��(���f6�m�w:͞�E
�[�l�`���dЋS1Z4�`��:�=y��i6Dt/�ۜ�ue�őg+���wLY�턀\]<���Ff�F�s���V��cJt�[��C��B҆5j�7_REHy�lbϼ�Yq�RM�KN'����'�.�j����h�E瘗�pU���֦%����^x	��u���aa�I����P5_\ۉ��W��*�Z������l�	�r���2�(��{	.��Êۈ��r%�s�.���f̙� �'N{\�y8�d�e�OVr껼����w.�k���:�1��R�.S`gP���~̺���%�(嵛�<ܢ�^������q,�=|���J�p�"�ʐP�<l�CߗA�Y��^��W+0M�� �6TB]Β���ُ+P_:�rh�x}ț��fa7%�+O�U�r?���z5��\lm Y�����`Ì2�vs;������1j�ܫ��l��;����������t�Ӛ�E!h�n���t1���Y�KH챃%z��2����У��B2 D�pxO�ށR�T�/���EkN{�KVI#�@Pˊ�n �=�0��<>�/��ҫ���چ	�CX����}"�.�8�O��ǕB��w	
�]S�����[E4^����ꞔ� j�o���t��D�w�''�ri�E���{�|�C!����C��	&��9�@�z�=G��c��r�f$�,� _�߱I�V���M#�e���"��qe���r*M�!� �Zύ���-h�h�>0����	���-��ͺe��.F?3��,jFSm�\D{g�yLO����"�L��` ��E0�G~�q!=$�0?��~�Y�nFf�u��<.��G��}jqO?��C�[ib�i\t���Fг������a!+,��Y߄'��yO��!��#?��G��,	�
���8�T���J��[w�X[.����پx�Ɏ�H����=�æ0�G]�Z�6ug�huTퟙ��τf���f�at�������+EX��dj'�a�~p1ȲW�Sn��I'~A��.c���7Q�2�gя|�!���i~��n�~Vbc��O?-nIi��4.���I���K����Y>,�,/B�X{�f�kڂWz���I[�3��O����k��3|�'�����$��((x;�Jȗ(X���(+ł�0���˭����E�J���y)6�o�q��}�D#M���k� 4U���gT���B�f��d��_��{Z�q�� ��X��fĊ�_�.M�"�lp=�� �K�*[u�f߫��F��
�8���R��@"����|*���D�;/n-�(��%��'1؅�.c,ٳYAT���u	4Y��=އ�"��br>�=߰����f�GA��k�|ɼ�+�v��\%�B�c�Eg�}$/�|%
z�i��'\�*��J��MI�DQ��^��D��4Y�`����q�[E���4Bϲ�]�aa1�/�|'X�g@�]����L��('�yK��ǈ�t�a#���^p�q�\��a?}�Zf��}�19�7l2˾$p���6C:=b������5��Eg�@��bQ�fЇ~џ�!fn�Ź��"�ߜ�/�G2����wh�B��3OZ�dP��ły����|��j.@��~k��C"-I$2jg�X~�a��K�{��O�?K��@���y�h��w���zЗ&8�xݡ�R�hy�iMG�C���n�7C�הCO� �U�[��4[�*�[�{��\o ��E[�l5��׷Q���4U�{�g��NB�v���_k��HvN� [+t�
�,cz`����X��-�|O�Fh� ��i�a� �FM���M"8��~E��k"3\L���Bө�l��4��$��E�~��lջ��Y��E^jG����Z��x\ ]�Vҙ�1M,?O�N�K�Ai�ݐA�A�����f�+��I8�<�'��TM��AKV)�ƳA����,F�p���_y�o��FJ>��y���h�J��X��� |�c����E�Xsu4/�D=6>����;I�meF���猅��#�����x��-'�_(�,��:L���X\>�h���-�*�ө]�"ى����V3gB�:�Tf���A��p�v2M���k���h�U��y+�p�]Q��<�*�!��w`,�W�(�]tHYI�R���Wqt��!)�O˕*�4����Z��W����$Fԙ�>�[����ۥ��,3h

������uzi�ޱ��7���8��X��b�(��8V��4�zo�۱�m�~.w8�3���9v�C���-�in�+@���X�WڅJhe��c,���J!��%Y|>��/��F�N�!'����C�}�T��Q�e���Z�s$q�F����*J_�y���'{@�yW�C&C���G�w:�K s��/84�u�sl�qVPd����j�����W��f��>EQ�3��1*������6��-�)�8��|�����e�^�c�KH��������U�y������Y�H�	a��^�Jz�F�ʢ� ��}J����{�Ǚ�Y9�7 �,�e8��~���b]���k������
�,r��P�TP���,�;����Pc
���jE�5w��.��-zqGp�����e}�,|���k�}kg
س��8����l��Of\a���q\j���Q�y��A�g"��to{�+`XE���4[�oኂ��X[�A䎕>�s;�e.��3��'��ϱc���R�>�f�Ԣ��U���\cl�3��P�j�)NB˽��1G������h�*!e��s��,V����涜+�]���̺<"\��y�j8 ���4W��6w;�Ysv�b��}�����]j��.t���q����Z4K����s[Y�)��"����G�� k;jt�v�'	���7�LfkPѩ ��m&AT*��i(��3?�P�o�SG;��v���㥪����дA%�ƃ��&Ѳ�
)����vH�F�w���Z~�7��j= ���y��f���&)���� ���^V��5�t�E ��9ϯ�Xw^�DX��kPy�z���C�\�|If��e����~>��8Iz����5�iM�s�'c%�빽��h��O���Z�-Z;�P�ߺ��d���|�i�S�$ =�M�5��, �*i
�.ϣ���/Xf�T�ҭ�p�j�c�K���+6���3=�X}�v.aŻhК1% �a*��cc����ZIy�]4	�l�����
�����W��W��G>sI��8\�>��4�7^3@+}H:���m��OO��!7	�c��'�i.���`E�7e�=B���gE��J޺�p�F�7���H-�H`H9�^���h�hg����nW��]�)p\�*�|u���.VT�l2����H�xF���͉�e����+]0K��k@�x7�P|^#YLwq,����Im��4�;�ӣ@����"��ʉ��+̋���f��r�\ ���H�Sµ�	@�2F�>?[����%��@@�?��@� Jq�������؜z���P���R�mX�>x35}��_��*,y���L!$^@)�p�7�� �[�ioa�$���^i�U*�_���]��et�&6i����NE�a�^��W�}d��AvEk����E�yi�L��1V����~Δ���s|b�e���=9�K!��w��hSц*�%Ö�}XAwbr�ބ{(�糡S�� ��]�e��P�n|�3�`I�i��wE���O0lkK�˅��Y�V��.��W� I�K��h�V�]ZľaN�VӒ��2�FB�@��f��6��γ�1�#9��Z �������YKO�g�}��'�b~vF�'��uB����b�*
�P{�8���Vc��:��9e���D� Pr����Q1)>Ql+�(�|�}�ƙVc�5�V?3�B\��Ǌ�8P�;1�E�=�r�x�=�>M�y�S�WiU���@n�r�0cn!q���bUy��/��@�6��a*܏^������
���2hL����=��e�+A���|����Z )���[ap�v�JϚ�T.Vs��UFKY�1�o*1��5�.�, ���)f�7����̙݀�1�/j:��#��\ֽ(��+�Ox�2O"�R���f�ڣ���y)t_Rj|�V�$��U���	N��E�'%ip������b��ŏ�9��HJ�Z�;*G���r@.��ɴ�M����Wo�lpDOm�;�����)��'ؠ����_��d�(!}q:�E��GɠX�as��z��{�pu+D�b?�������g��Sm��uf�3Ur�j!1"��S����� ��d?VA	ݙ��z����0iH�5���t�<��t	�*����y�#���dYS�I�����G9������$�8Ȫ3{�o�`3L���\�� ���%͡eK�ϡx.�k�z��:��~���u2����V��"����Cݯ '�n����اY�~��(�+�VTY C$�W&'��)f��g7��O��aȶ��UI���י��o}
7����q�^g{��yp�s-홐�0��WW�Jts�`�Ĩ�C�
�����L�"b�H��`�4�
��T4�*�_��4�Q����y�ن��:8ǰ{e���b�&����k�c̏���XK����Ǜ,�gur����=�=�/������1��S�[|���O�hz����?{�p���䊆�3
�&*����!�����@�ߧJ��j
���D��9��lScbi3�������di؅��ܹ��-�ףs�V��΋([}��A
��;:|5:/vy�.�@�-z��3�߬r����,!��vJ1�m�Ug9�����H��l`TB�}�)0��bgAf5�D??���$�I�^��o���:�0W����J	˴A���]5nj��a�1Ff�61���5��#��;
E9kG�+)�
>��Z���A1�}b(�Y*�o��]'��)�k��k� ���0^�S��S}��h��n*pm�f! ��
:{��C%p�-�
���m7�Ft�G��S�¯��tR�l��d��Y�:�n4�@��2�\��ZL��xgB����V�IW�S�	&�m"�t�K1�t&��J����r� �7g��u��I�����i9I�f��pz;vSP��ȿ�v�Ծܽ��=�u�-��:g����9��Ax���-Xg(�_py�0fe�E�Kn����mro�bE
8G�:*2���_�_��[KjE�?2�81f�F�(=[���.�y�����`�φQ��ɾ� ����Ԋ�HJM l�S����l��fv-�������6�&���E�e�1��Vm!Ю��}�t�S�X�W	}5�����eD�C�d�p��;ѾF�<��;|.[[&X� ��͠Ak�F�ƗkK?pA&b�������{�ұ�+�v��T]`���#e @�cə��Q�)N���ϫJ8֗�!�-t��[�ES_��;��ʃ`���0�NU1=w1�ѻ+TzS��S^X����Y?�+���ڬ���G�
{�G��0�@���2}�o�6�X�;��'�gf�ɪA�c��|�.;��r���ӄ`	�5���^��՟��GO��ԚƦE�I3�E�m�-�Tx�PhU���Y�`����Qy��{T�-��|�>Z��"�UE)J�N�sVVŮ��f��j�J�{��O�p�yE�R����4���?ْЮc�Z��D9�iWt~}B-�2�onM���._��@Ο�}V+���)C]�� ��r1�xu 8��1�&�ʇup`�;k�+ܹ�<�.1��5���R�ȣ�O2�4�M{�A^���>�d��Jn�u7Z��,�� F��_Ww�nߕk��{�����������')�7�˲%������;rט�.@�>�`��"��R�[G�ůr�9ﯯJ,"O�V��	Civ�E�/�NdL/���KH $g���V�[���9�`�),�9~�P�%}��#R�v���с�T
�/%H04�h������!�?�/'�Xk�~�����(�nD�$IlŨ�o�����YdQ.�p�,<d;�6P�B{�Y��V��u��k�]%�A)�`�+��
�nKK�n~�kAd��s�E�Q��\z������~�r��y�Q��M���i�H{ɻxtHa[�]oB�޹W�'J^2�޽���3AI��ղ���|K���v���\�ze�O�>	���6���YR�Ȏ���i_0-���Ԟnľ0����}�n����t<�Ġ��͜�r�
fʈ[���
�+�t�*Y��x��厀Z)nwL�Z�K/���,<2~�:���]�lEF'g�D|�&)��T����.]tU������	�%�Dd��,Ͷ�%�T!u��yL�Ո�d�jT�)�%`��0��x�Ȭ9Oٚ;�\��� pK���4s�l�(yfA=��"��z�^?RM����zY��H$�y8��G��U)2"i�n�%M��:̝�}���v����ѝ�i`�ߗa�������t|�v��g��� ��[79�Ѹ@�_`���߰�-f@}��˜�s���\��˼PJѩ�UM��$v�������*oLX�nP6+(.g�C](�v)3λu��o�or���bN_��B-���".҅���{?����.��2�.�3Oȃ���ZG���P�>� 2��+��D�V/%1"Q�~�ʣ)�V�E�II��K�xzsD�@��LF���'5V@V�dV�-�!��/1��)mh�V76Z	�g�c�QV�"Ėu�d)|�-ře�LEwv{P.KV�̵�|+�&u�A}��n�f��)�#x���	�&�O�<-�V�`�J�Fj_sdI
r?���L��cnA�S��U��s��|M�C��a�N���4#��p��-	c�6@R#�4��P��f�eϋ񗤍 �t�8�6�I�O�7�����)6��A�z�hrq��VB�Ӱ�T�v����?��˸9E��sP�pɬA܂���%��o&.�������%c5�\<X�F������ޚ[�V�Pw|��K#����)k,K��r�1Ǎz'@� r��\��8/1<��[��JV�S�ԁ$��}�P׼�)�SL�"/��°��[�~�SM�y����0��G���Ͷ2m�|NXE����Y׀k�zUi|�b\F��A/�Ēs���M�#+d��b�(q��W�E�@a�'�Y=a
�����4i�'�s��h�X����⋬b�V����(�1� �5��u�B��>ߟ{���jne�"�~"R ��"��r4ٿ�+g��h�T�W�Ee@���i�-g',��Ui��So�Q����Qu���ԃ��fH6C�]Y}_�ꨩmB��8+��|3rr�����za�t��WB
�2�t�� �GM��W�'"O;�'u�5��T�#D�p��tU��T`�)��S�9�R������ǵ�T����a�l,<IG���>U�#��͠> k��7w��%��;�vX8hU��[�i!�Ӷe�kM�F���񱇡�+�א�x~<�zϼ3��(���3���(ЊK/#�jZL��Ue��I��C���U��Տ-���[ B���e�l�3R ��9�ɾ�O�
�O:�D��G.j'b��ގ�x'�	�m��+���T4��|��8�v$�e��n�)��AFd���A��P��4Di?wq����g��6"��c&�e
K��،��y�J�?:�`G$I�X.Őn�C���(�$�/�i�*|P��]JʒYQ)`9~���x��kh$oˮ|7\=�j5�����pf!髇���l֍���ے�؝�V����������R��%#�#��;���	a��B}�\�3���L����x�,�_��Tr�t�^�=lq&c/��n\�͈�M.�|����b ���a�~G\�hCC��-�>���B1��lr��������S����׸�uz��z@TLc��~d��4D�Bգ_��[�� �NM2Q��^���I��Q�轧)
ZbL�}��B9;�=�|UG_n?)�������2�[ �i�׮x{�AL�w�u� ��`�
���%z�Kw�?�b��0��nv�Ą�~~G���}6U���@xbX~(v++�$R
"����Z���fd���Z�ͻ.Ҁ�M�`8S��Q1F<��s���*1E�0�����D�w�b�D��r�r5��w��.Qၻ�k��j���$˳P����3Y�[�%7�� �{��S2��/�[�Ep,�Fa ���=��i]p#pe�����6
D�VO�� t��,4(>�n&ַ�Pd��[��d�yj,����(�@PÉF�vσ��-!q	����#��e���pH�5���k��Ǻ��-G��f��u
�}.<{n�22��Ҩ�%!NT�#dX�gv'���4���`4���'O5�qJ�%7��m����8Gk*�j�#�u�k��Wx<�s��� 7S+��"��kM.Sim��8J�����{� 7z5�u �U9u�`}�\�U�/�cU�e����+��{_.���{mdi"��I1``�p	&�{�|� ������ �%�A��L�z�/��@�M>CO�km�'�H�Ƨ�Վ6-����z�Ŧ13�0)��Y�%��`A�:e�8�������k�6Q�O��5�/ �b�A�W�K����An����70:3�p�s �-�
�f4�S�>�7S4iSL�8��w�~?�Q�1�����wk^a��IW��|���&���~,���z*>$׹�8��'��b��u6ֹ}���Tf����ogbge@��$o�2_���E�+�QX��\�m����͚����dg3yUt��26�����o��[_�H4��b�夝�v1���3��U�zFn��a����h��]Ig���ϭ[I�u	����>`X��65�n��%!F�m��" �>��%�	�w}���E*P ��'v�O,��e�f"׵;�}�o�� �Ŏʿ>��q�!�a��l���{U�$���RV4�AE)Z#^k�f���ngLU�'{a��<����'���mb�Xb��R��@��V�[����L�=n��r4��b��Ӥ!深��:]�azp��8����R�U~�4zO�����Qc��Z��>��E���bv�&��ѻ1^�`�x����� �޵4���B��fJ�@�
�@�Ni�C�ӋL(�?f�x��#泇KjұhnN�h�m��z��k�/�seb��f}���?�$F��y h$$��� ���&Nz ~<����+(r}a�t����j7�&�_*KK(��Y�_�߱��%-�^Q�%�E"f3�
؟A,x�XĦR�w��/b��l���c+'��W8�F�n��;��Pó6A c"��N�����%��ơ� DB�Y���ڀ�ĮϽ{��,6-Vcp�ޘ���'�p��\���xdȥ��n/�(��g0m�` '؛�!�Q�:� �3�]�4��~PaS��J�'O�(L��6I��]#p��%��l����F;ъ��w���f�EB�Su���9=4�l��C%�����Q�1���!��sF-r�*���O#��I�}�Z���7�R�Φ�=Ɛ��|f�J<5Lw�B؉�U�`M<��PW怛��2�_@]��Ļn,Q���3LƢ�[[P�Mۃ"]�f��a;A�=�>��݇�}m�6���ả�=-�Q��!#�V�QI!kY�40nO��fJn>@Y�<C9�{��Ws�-ގ@���֫6��6?l)	|.���کc���6�W@!�6g@ђ�Ԃ���� ^��M��㊈-Z#LIǤ���h���Ǯ��cɬ<P��0��A`Z��M��3G8�'���%��tP�|\�����e�@���/����KⳢcR��[������B�t�L��ˠ��f�U�o� �Z�ԛ�U�e�
0���:�<|�h���u%���+}�^�S����L@��|��R�+�#"-��}�g��M��]�Sf���È_��=Ϝͳ�:؋^��U��:FW��_V-���#�R&�
5�L�5[���zuh;����±�;�^?&c��xj�M]�蝛"�����a���$1]���yu˲
z�04̏o��d!Y���O��3���j��'�x�������	9�C]�m��Ck�����������Ϣgk��/`��[�B�ɒ�s�1P�2�2���(h�w7f*��F�{ł�:IBѶ+��/��8��0�t��c"��9G�	��7�-_�V��|H(V|P��"��2Ϫ�A����&?t= v$H/M���b� ʃ<��>!���m���WP[a	� o+��J��x�Y@�]1.�-��r+��G�PV3�o�:��U��������ĳN�'�,�U���H4:b�RO-Κ�r����+�OX�\�)��vq��m�#.�.��^K�;.u��p��*C d���d�j�V�X����b��S ��lxs��N\ۋWf�Uh��,b��Wj^i�IzjDs,����4�Х�`jN�K�]E˔�F,iy�ќsY������U��x:���!Uי���Е�MX� ����IX��U�y���Q��.m����VײB5?��d��"�{
0�P��ɿn+l��>1r�"�ݎi��I4v���:�HA��pZ๦�HX� Q�qA����;j���ɃT�f-1��i2ꑑ7I6��s%��By'A�����&�$�}���m�
�����'H�en�;�7����>C��V�X�\zF�1ى�p��!gү&Mp����Oٸ��v.�JN2�-e#\aʖ\e���^6�5{�Js3����3	��[�+��(Y�M��z� =�4��4*����x��*#�u)®l�h0���M0hτ���ceESFc�W�C�	-�^��Nd��᢯�T��Ú6v��{�tm'��<ͬ�Qx����_.���K�&�M0O���7uW���@=��n�Ϫ�B3��1���	����I#.�\�l�����W�^٠���٣�Lo�(Y�p{N9�R7Gz�n3����t]��B��{Au.?�h�4,��h�:mF?0v��#�BG�VFs4Q���)e�ǲ�b��d��Ls��z��hgZ����8����,�΋Ь�k���! �L���e�	4-��,>_���d�޽L}�4�$� Zl%y��dVsH�u^`�#jy���?U�g�Ǖ��r���������閕!���s�ȠU>W���<.��Y'�gv9���e��*���C�'K�����l��뱆�G�a��c)�c��/94�ajSQ�g�H4a��qA�T&�(�~�9��[�/�t���V��fE������E�vI��_�	A�?*{�i"�i7]"%�	�d��ʌ�;^������������$��]d��n���h]Xe�)M�lK2��:7���rn�j�`kC�&7�R�ߓQP �
�&x�-���;�K��_���.H�U����@@e\Q�7�x�覆�0ca���	�N�6G2�Պ��(/梥H�t���<ڃGHZK3�'��0p�e��(�:���_��T�A&�����_�NƮ��_?�����(�S`V1�l��|G��҃���g#r�!��~�1�w.Ũ1١����"b�Z��:��j��c��]rM�%>�hmo���	yX��aqaח���>�ˑ��+�	~�b���l�wU��9*F;�䙉�B4��5zh<I��g|U�C��ږ��@�m�`��m��;�♒ 5ǟ�޺�Ǔ��en��i��n�H�y�}��1����E�a�<�Q���#/Db�T�X�x�Ї���d�"4��h�a8a���t�V��9��o\Œ���p��y�ߊ�>@��PA�g��X�PW�����:�]<b�0Мǥ%�*�F+pE��|�yI��*"��^�4y˨Tr�2�:6�Aÿ����1��V��P��M��1,3�4-*~�%M�n�R_u��5����	����']� W�n��V];C�(>�kP�߅�G`�I@��vF�`>!��7^w5��F�~F��9+������q�����I���[5���'��jF�� �k�A����W��oia��곿}j�B���ab�Tc������Py3'���̈́�>r�ER��igq8��*���l	�����}�*�h�+(������t�>c��g�}k��ɹ�������¨a�T����s~QI��cy#��S1o[u���čp^��r�gr�$BW�-���v�[xE#�}N�*�h-�D�[r�s��4�V���j+QM���9
���B�"K�)��i�f-���^�w��fS]�dhI�\ -�\~^d��|����0j.��J9�&|ձ-���x<��v �$����_g'�Ђ���ǧ$Z�	�$ϦX�J���2�;0|>��˒��X��|�r�C�)и`u|s�y����-Q�Y�z�]��B�B�7� ERfF{{��m���N�:O�m͈��Iu;ZX{�pv䤻=k�G�[��[Ӷӱl��T+��ʮ6��V��L�N��ȫT@j�.�0���4G���ÒMk�{�*ii%q��+�Wj����Z�P1;D�'��A�d��07"R �x�ֈ����&�LP����>�č#�^t�Q8UR?j���M���"����� �PH\�h���B��̿�̚�0eS��w��ȷ^��o�"Mu�_�R0�K���q �o��k4rL��]�+��<qT�n<�w�CI0N�_�}^_�H�+羽˖P!ߝ$:x�٢u\t���~�����s��"8g�<���ݎ!�cM�3�W��P<C�SQ����H��H������ne�s<kQ�7�4XkK#�jl�����2���&�
�h8�ӟY�51�;�<��*�ɉ��,V���(�#TJ c/=�`�&[�v���]�a��L7F5��#ߚh�	q���}��2��w�iex�3?��sZ��]L�Lֵ�{_5�,�3�9.AK��עn�g��.����KJĪc����)(��Q��H5���j��D<���LUs
��-M�.H$��?|Q�(r*%`$H�\y�W�7�wW�2Z��a|�W��	��-��,���l�ԩ�4�3�^o�歞a^���5�vs��$.�+_ �NE]�:�D�tSgޝ����/ �!�����O�Cce2�ZpQ�+�$�O���Z�
� _]����W�7X�N��h>\O'KN��3N"�	��Jt@��p�4���5�j�Ja��}��p�B�0bg�sr.p>�8��Y>��Ƞ�(�c+�*w�Q�U�Z`�P���v��qAB%��E�ϓD���55E74����*b��sdm^��[!�����)٪[LI�~PbK��8c�9h��DJ٪ĭ9`��C�� ҍ�\/�s{o[8V�-���n����29`UػBl�ƥU�6��gWv���Q$���\A7��Hk��oQ�6T�|��Z�D)�`��K��|j�#���K��ta��2��0���7��ȭюl"����=�|��K�utۃ��i�����Bt�!�u=`�{|���� 0$�V/$��Y�I���k/<�%��&Lg�<oe,>�����o�v�m����;�c�l��踐'f�KCX.v!y���]��Q�������?�3.�.ݱ]y�i;�<�X���b(��K.�⸂K�$ͼ�Ts��3,��L�3�����X��a��+�J��Cfۿ������ ^�^p6����G�����gëMT	~����䕍ݪ�]�"	�1P�X��N�ׂע
K��I�v���8@��\+�M�h���N�D�Ϻ�4�9�j��@�m⡥*d�-���#�YJ�-}D�!Z����׫�T��%���~@�|z�&��� "���fa��՗W�m���� ���E�H/�vJ����ј���Ӝ �#c��IS̍������D	�ŭ,U�Z�b��(o)h1#�^��n`fO�I���ʤFR'�8*ΐ�c���j�� 3ۙf]����L,*)>��\���V�d�	���V��B�R�A�^ZJ�ԛ<{�!��:jL�z��``Y?>lK�� {�fR)']�Q���x����GW��SI��7��Ymt1K�!��ԫ�E���X��� ���O�[a檳D�,�,[�(%-�+T)4��f�duɅ�K:�2�t�����@>�D�Ր���ʀ�T$�=ԕ��8mjL�>�����C2hK���ʚn���(�T��5T��U8:�k1�/�+N�����M�: Q��9 �tu>ut_�-#�wD��S�ǩ��ͬ�j�~��!�Qp�9��Hڇ��O.���|�FB� �u��^VM&ڄ�_g6Ǻ$"��P�Jb㚔kqf	�s�ٵ�0t���YFl�qxb��o�aY ��d}�gs���F��XS�-�H䒁���Б[D�ժ�,�3daQ��N0Fjsy�M��f�04?����(M�$X�?�R$��^�և�X�_�����[aA�a���o֦6��]�!F ����������:��~&�uz,��p��RJ���;��@����C��Z_�1�Q�<�mh_A��O��!wc�y�4�!���<Dc��F���Q>�@���>��~j���^'�
�����V92	�

�Wj��nj�RU��]�@��eC�T�e�-��l%� A��n6� �t�Q�z�$��=2.џ�M�z�	%E�V��X�.�����/4�ݭ�\��]bC��$;%�*%��%u�P�)�ө�<R���Ѯ�~��xAK"-�����ۺ�{�j��e����Kg%�3AM��I������j�r�ڏ3ab�.d�����2_PT���L;.��l�(bO�*9h7�t�	�g��2��~���6����+�͏DB�!2��:i�.��������(��z�����)�T
@�� �]dF����7��"��4��Ӕ6$���L�
R���5n��2	Lj���FB/�����U�����CՈG�K�6t�3���~Qj�n�=ޏ�+ڕ�i�W�{̍ ��U�r��I��.�x+�Ղ/��x��p}G��d>7�7�Z8sU�S�ڠ��.)���F�1y��R�_S��nd&������E��7���y�������r`��-)`����y䴂0��7ˮ��at���d�	릓�ҭ|x��)�Z�M�>�NE(m�ۦC�5ߪ�ʒ����B,4����!;������&F��Yⲭ��[��p����~���Ϫ�w_�	�࿴��y��'�/5�������@^	����|Y-:���CZ�հ>#zs�\�׷6�V�_|Br�֕�/aD"D|�I�'Ca����$��]�T#����{:C��@Xf�������͎,�/Mi.1��_@7����c=�&|_F T�j�̊����3���������@P+vgH6=#���'ǙCO�sW-�&�y��V��A�_瓌��+Za#��YТ◉��?Iâ�a�.�w�Qj�
����sw����V�_ hnК܍��y��{�KR�O����.�=KE���)���}��e<�/�jnd��N���#��I�j��fR�YQG��ʌM^à��#FJ� Z��#���̞��k��t�n#��?V�.�(�E=�W&�����h�<OU�ݛ�8�0�,M��nNo��Af~A�	c!��ۄ?��&����92c	�.�b��U(�+T�?�Ω��LIզ�^J����gL���.؎�JhN#S>�R�N�@\��z�ٮ2�P鍭����4�(�ܯ�db��a���̗���܏*�`,eDj�N���L��FlP�9���{���^*�����kb�2��5v5�0A��--c%w�eq	��E����I0����*7�R���N <[z�u���$������о��و��2w�f�rW�C�ìH�w�q;]#��K��ˠ��Ι�@�Ü0����ה�m>�#y���i|���y:o�[ܯ?�����5�{9P�/!�D�)�6Ѝ�6O�g�xPd�,�ti�[�&�ٕ�갗�R%��Ώ������b�b��χ�����`Ղ� IVT�Ԗ��Q޾�I�A+
%�!^��2��Ly˳_�!�.� ))���ʉ���s#�~~C^G���h�� z��-Y�6Ui�ם��)�a��sl��~�	�-���ჾ5�A���a���(ɄUJCs�S%���:f�5O{��?i7�:��ꕨ@���]��xA�*��+��O4cK�
�)�[{*�p��ԃy�qۓ�r�Ͳk7v|����a�Fд�S	@���)��u�6H�fJ�1��l�2G����}8r��򾱽��"��Rhr���?��j��Z��UbhIAA�9�0�&};N��TL�����ezaGDI=���@�[�p���݆��MV�]{�vn���@��R/���&-�Ųz�Χ�g��g����g.RՍו���p��qyfR�gЄ���I��.Ys��u?]�������MW����EAk'��uW�]22�6���Nhe�a(U��|����&iH^>嵻�˜�#���wA	�8�v�d�laް�K�>7��><�΅'<2�|�Ѧ��4]��`�S9��%r��\c�Pt�1�=cr��/ݾ=�
Ͽ�2���<3���zo�E,cc��"$����+�BVQd�Tf�����֢	@��pj!�V{�χ����٢-Xr�YϦEV�G� �c��;,%��l����m��k�<y��*U����=�d�z���U�*Y�o��L#O��U�(hIey����#,Z���?�2�AG��R��[��i���cpuETu42��� R��	�6�_��[���\��}p��n����%�kq �V�vܬ#+�?�/0'4�N��`�,0��/c�[o/�l�'
�:&�����l�O�?���*8���S݆���[�镡�Ǝ���S̚c�kq3��g=P�؀������η��#�u�� g:�����~�qO�A3�RR����� c����d��X��#��ᙲC�i��R���>�e2�'������Ń0u@�P�2��L���d�pw�{Oc��AdJ��jO>վW��O����g(R���nֳy��X/-���+�1��U].�i$�=xO1�����sH����٦^~:ކ�(�.#�k�ǇC,U��`^��r�� �P�1d�XΣH��؝��z�`�>��Cn�3(
k��8���Y�̋}�x�,�Z/y|�~|�i N��t�w���ݚ�"����c`���$�PqTYU�9�x���/��;���� N����x�� ���*q����o=:`�#�7h&p@0~���_����R]��n!eV�pʮ>��ur�$vy�'qG۽���ݶ�Y�qѮ�hg;�A/lj���suŪ�]���zhP�1W Vo��?��hɪ�[�(�B.JN1�m4�X��6"X0�����,�|8�7|1����@���E|�Eg�����
i�c�a<�a[$j�������`ђ��k��|�g�V:S'�,�N�_��"M;���j���9�!˅�U;�)�b�o�YR��:62 �x��7Y��f�wJ}fU�����;f��'�N��x�ǈ�*����9�f4�F*�����|�f�r�iO��.:R�1/�)P����U]��?��#�.�~ė.T7ꖻG��K�x<���Y�}d�*��xT�)S�BN.��J����c` ��`�x�����
0��.mn�p�"�7+&!��VĻ$���4j���q�txOJy�Fo�`�������Y"�`J�Љ��r�L��d�#o�����gCZ����~Y�|k�>0)%*��ζ6��ѩ����|vӓ�&U� Zu��y�ݍN�N����z�d�{)���!w5��+3���p��2�g��:2_O�G${�ڴ�n�s�%{�|m9 ��r&w���tH�+��U����dI�<� ������o:0�J��wpg�)H(�rW#�g?l���į���&Ͳt�W<�5J�_]A2�U�!�I�#Z����(-g���HS5���b�[H�s�32�#Fq�L�~�t�@:��^_�eB?R�i/��K�c`��BiqUJ����oOɦ`���h�J�|V,���lv�����ϡ��Xe���N��R{|�)���L{=�=�a�F�t�CZp�L8%�n���|�l �m���&�cB�pf#gT��͢4VM�a����|��vΎ�X�!�F;��@kx�Y��7�$`K�o{�-6+��G�@2v�ٌ{4���*�|9k?ৃ�W7��O(�;L�V�w�b���b%[�r����"o��Jxar��2��%Dg�X�׶������@��J�ɫ�ͷ������b�E���wi`ӾQ3��j�RqXP�x��&T~�k��کNl�Z)�o������K(��R���g�?�N����E>��w���c����{�Z�����e����z�\�Q�}���LyK�"���͘8�xs��y���+��l�W����/}�4���-S0k3���0������ټd�[�;�naEYi|��2ZZn^��%��:�	�:��@�f2-��ʵk�:��w�U> �'Z�X2�L���*t�roh�w�Me���~c҆0­ ��
��Ճ��,Oh���%��r�h���̖,d�����X��I�o�� ��бK����.W��oj��Q�|�����)Yc���N���M����s�Š`�C�h}}/1�ɽ⦙h'Nib���
�u��V�VR�snj����?W����{�Ny�{��ƪ��]��Շ�n�Q��q���3A���`<ki���^�Z�t�`$�p�ԡ��{i�$����_��̕~��b�'�I�À�ף)�j%��A�ҞX)��x2�7=/;P�	rԃ0���8�D� yW\������W����f<� �z@n����&J:sp*L.Ie�E�XO��} Xw�y��$��'K��g�-����Xn�7v:)]h��cNV��d����,̾3W�ـ [�2l�t��e�$�C�M����vP��x%�0�/S�Nd�X�F�&ݷ;�(g���s�SF���q�-(�]�'�џk�-�Q�N�< |�#,��Re�~j!��`��`m�0֘��ef骁��N��i/���GF��]�c�P�)���U���%��u��U�^3����P��$�E���X�W(E�Mxty�T��S��m�Ӽ�`�IH}X�����^�����>��N�ugz���!�/�Xu�P��iu8bQ��P(kJu7�h3�7_�q��cP�Q�����:�q���aY��@�í�q�Ք�M��)X�S���:k����>r6����8�R�+��q�a�W*Q�qf��kW�5�.�a�\{���[��]�KD�������	W�̾V�<��0�o�֊A΅G�7SX���	8��ǘ�jD(�B�\��/�w�xW��3Te0x�Qj���1ϣ��������61�F`kw���ݫ�_g��g�[o��E|a��J�4+�Z�apq��ז��m�[���"2p�3#�$9������Evp���-A��!2d�����t��#���3%d��}6��5�z�
39��+AT�Ad�?�BQ�&}����̵b��֍�� ���X���/�4�v�o3n���lj�y�V�s�R�D��@�r���ɟ��'�i>S�L��:��`�Z�杤�+k H��"�O���@b~�K�ˇ|1�e�Fq[� ��jad��-��ͦ��,�>�ljU�!�-���GK]�Ҽ5�Ư���ä����+�{^�Tȥk�X����y-2�r��!����?w%ﷵ��x�ufy�#]��z�%4`�<K��k��v2R��2@u��pJ�܁�eC����iJڠOʊ}H��`ڵ^���2"󸀾�@qƶ�ϸ��ACF�{ ��	�\�J�d$�ZR	Ѡ8v��q��y�0���CNYb���J*�\mw���=K ҹe5�(8��0�>.|��bm����b	@,�	�G�	�f>�E޽��Z��0�J��3��ɺT>�9��5d���&�я�M�VT�
:�%Ӑ|b6x妈
^���ą �=�J�P�i��l�svk1�U0t�^_�������j�T#=���O����HL����05�L[��A���W6���C_~J�b�uۘ�f0�ߩg�qy�Ǻ�����nc�֥M���@�DDn�2��̱��u)F=Ȧ2��^F�����Wu�ȕ�O���)�4�2��_�nT�e`�<�
���t�qT �^[v��Q)��N�:�4�H����Ĳ���JJ��\�HٯQ3޼��2;QfM��R�ݨ�	��n1vI��U����&M�ט�Ї:/s�L�ܱr#{Ƚ�D?�8�<�}<&u���U��k���?։�͚�4����6��^�Lq����8�Ez&��&_y��c�ЛI����!�Y��3�К+��ݖj5����$th1��:p��	��;D&���R��4�+���gk�fp�8�i7W�����.�����UB�N9Uj�&�pC�Kch:;n ��i�����	v�<[�E�bߧC��wh\r|Ú�W���� ����[����|�&_ڋb�K�1���v��"p1�+��n�"*����ϊ�8�r=[�4xZa��]�|(K8�NV�1�˶KQ|���©�Q�}����c��Q|!��uÝ����9���f.n�=�Ğ:�ns�}�AJ�)��u�})7|9��4_7����dծ�*�B���"R�W	�����UD!��3q��P�@�g[�j~CxKZ��2sB?�h��c������QM���mf_I۶��9��!m�:!8�{|�V��h�W��I����/#��-��d<~��o���UB�����l���<���������H�����!����	��7��42�d�;+�91^��T�>�1p�ܩ5���o�uP��T����y	�NY�}R���C�2ɀ+�v�k�$�si<�}��S�h���ʓ�J������)���"9e����1ZUd|�`���C�70��J��u�Ш��6L�L��^W�+��V��c�y��(=�X6�x�"|�ɧŲ��3�n9��������e�[bf�2��3�(�8.O\�LQ��E���
Qh]V��ʽ<�L�JĮ�u攨�X6#�L���a�kcXQ�i�h0*̝��)�/��!�+��}�.���#K��u��	�n��gL��btzS�~�|PE�94x��lX-�џ�x
ʿ�m��Bn1���V]'����o��xn��M����ƙ��tP�5�v�O-�岔�.f<��"N�"���ʯX8��l3OK��vE,�l��34��B(��Qsol����A3�z���[�9o�J�������j�3�79%Ő�;�@����S�V�3�S�V)qf(hݽ�,����!�~ ��:F���~e@8���h��sK���O�C\k�(՞7���H���L*�?L��>�?�Cͺ�q�g��Ze6c�3����nⲶ��k�Q�ꆔT�?��%���{��v9n��"��d�vP*!@�Xv�3��ۆ�M��Ұ櫪��#v-��7@FG��i���Zq��i��>��Ϙ�9��+�� �HѰ���ywe��T�&�/���11�'��O9.�Ld�Ҳ2��P�6ǝ�t^�����I�Z�Bj�t<���5D���b��#R�e0-Q@?��{��N�P�]�o���Q]���m�N#L��.��<�s`?��~ڼ�<->`������o��%��ҮQ`�=HUOf��T�U;L����qj���P�%n��?����g�ܩ:s�G�s0�MϨ���B6g_DS��ԋ�k�W��4m���a�q���S\���N����"T���xG-�Ē7]��4�3�Gp�Ӊ���o����%}܄��a8B�Ƀ�"U�� 4���׺�?��EV��O�����q+�Q #�nU�E>A:y휛��|i�}�C9/g�����щm)E�}�v֏�#�FD�*ܳ��lΠ(�s�.@���F&sN�h����"���e(��ד���g�=�����Ͼ�R�=hԟ)<,�����J�uM��9���֤/������(�'̜�f�w�!7�j��ihĻ/M�����q���uwЖ)��ē�ʩ# >��ŪJ��4�i�p�F��7XvG�wdJ�j�Iӳ+-�?�L7F{��f��� ���'�����]��~�BX1W���Y�i�b���]�voߚ.��5���Q��R��E�/��xs���'��<�gz;KӋ4[���$��N�R�s�P��1������)��Zj��z��x��>��Y��6@�\U�]�c�P_�t�F�<w[zuD\wE?�6�xV���^�I3Uz/jJ�Q�Pc�9����׫t	��xj�r��� F��� �PZ!y�IDC�얢�1NL9'qp���S3`��ʗ����~��S���i탼T�����u�a�.�<�$9u��i�{6���Q�<'�H���h=׬�|�4�40��2Y�����5i`�4g�Q��n��(�LW��d�n2�z~��P��U��1 �ec�{#�����6�߀
~輞���$���������Y���0�l��6��O/hغj4j�Y��l1�D΃L��[�ؔ�� �)ʮ�)�(��ܟ��ժ|f�~�$�����Rf��c(bͺ�=q�?n����U��o��b�/�y�N{��%{˾i���~}��a��e����E�Џbȅ뻰���:B*|�����n;/'w5}}gM�8�� ,��$���_� �hcE�š�}��K�Y��)۰�P���q���$߅��2)�
��ΆJ&�Ӛ�d��������A�tpKW���́�c�%�� �v��v���}���ÄD�F�}���6��@cﻫO!�I�xfk�qɊ���E��K>J6v��5�}�'�0Ѥ�P><���a�v�f���7{ڮI��A�ݬJ9�[��h��]�tE�v븘O��#���jc"��w0����-��>B4�),��Y	ۖ�;������O��+%}%q~�d�>3���`OC����'U[s���~f���ƶ�k��Ɓ�qmt�zl�'��� V>\K�w���y�����H�D��M��q��~��g]3)MG�ї6�*4�Mܖ�DV�-	6`� �+�J�&`Cv�i��T�H"������M�3�F�׫���JXLiGƃY�[D�������P>i,e~h|m'W�7KC������L�ޮ2³���ƹ(┶PzD,�����2^�W��CE�(G���� D�J�D�!5��i5�e3.����	D@���F"�c�Zm�<��,bi�T�r��N_ї��WecZ�+ةwD	�,dY:
<3}��y$�I����+�.,0*\��N:Z��)���O�#�u ��QĜ�������	W���K���8�-�X΍�$J��>�Ҭ���֌WfvE���^:
bIuI.������-@tb�%�dl�7�E#�wo|@v%QBT����!Ꟙ������(f�i��uy;>��T5�X���,'��<�)$[!݈�3� %�4�jHOaPЯ3���q��
��u`�a�֛V�@����ï-��N���hq��y����`TB�0[�݁��ZL����Fs���}a�oz:#RjΈ&���>��Bc�ƀD��G�I���[�n��F_쩈z�{&�)�}Ra/����ID����E%%bMV��κDKj�߰�?*�CP*r ���*�����.�Sǉ\
.��S�	;�tc�'=DF'�d�XF�	0���ꌉ����݄޸F�mP�iCLME�Ϋ���	�J���!S��3�)W���G�~�ai-DZ|��#+�a�}��0�"{,�����#�ܑi�h���<��A��_ʈ�I���@U�i��?nH$��*���4��O�}�k�֓ gyR�*T�����4���o�f*)��1�b	�)���l�v����ܓԐA���ڎC3�k{g0�"���
G�~�9��k�qo��*"��:8:���� @x3�2G�|_ȍ/���!�]�˙شnop�x["�BD<ɶ������t���E,�w���������H��� �D�w�P8S�'��Ɩ2�{xh��|�U�*";��Fb;��[*����l�kN��a�qR�9��pŪĕ��?g %��3ڕ�`D����k9�~;NN/σ�/eCl�֯2����P�{�9�X�5ىܴzTw�09�q���D[