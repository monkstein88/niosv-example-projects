// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
knZzWwZOdsKGkEht4am+7hJslXeAKhiKs4glHhE+RpgyHJuk5lB+WsxA3Nn2W4Gh8K7tzu0F3bua
FMRFBli7G/7ahN+NTFst/EKxxz9YH2z8W9Fvp/5PNpEDvq3nm5bdb/00tz1mn+Qf6mb2jvj/v3l4
eD6NbXKaNzglvILGIns1bY9r2C8W5V2uXfHV+HAONRZJeIQ1NLMaqlNcMFMDHrs4m7s5QSGZi4qU
Pb5OTerUZH1lyMa0kb2FlfnTxMm02ZiOhm+dJh+4X2PeCSJknidwGDDVvl/YBCHLiiRnqCkRv2d6
IHEXoWF1QT4lGtR7gX0wnDM1WP/JKIkJIj+cYA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5552)
jPD9UvKFlD6Lmosp6nD7prN0qitPd3OCgocI+IGZ53xHMgeIa6hBQamBwKImNp5z8/EPHBVhm290
gSYw+r3K3IiBVfGNvPykaDTqaTEWqk92dxZPxRPjKuFnoSHy8o6AgF6RZZ3eyBHoC5cZ8NifF0wF
8KRVcF9bL66JjV9Z/wgntWBRlpS0cXiiyadg0Dwi5zKLKqrk3vQE1uAFliy9e9uDBeyayzBYRGEh
IklaL2yBWxDBZY3uYoAKrgGBwdvLyLgt+MsJtulKedP75xgaowGxs3FGKDVP8b3mSdVSVJadxSaZ
BF7iy6b+RjYfjro1G6hW+Fn52JPYn+kgmwVcRimZ4ulnQogIgMnbKDYhtATU/pT9jHRv+X6/n4rw
UvcJCCNmMQlFOQXyzgiT+3J9zpQj4Mky+MTt/qtlu0s+ALvsBt83u0gNEGMBpmJbVA8D+fowliDt
EBBLrZHabF+j/ZjZgtCKUZC15Rp85dRmi/Zoq7qcgx/6gNQKn3U7DHZodS87gKO7mlTJOPNNVvYw
eXAGiSigAF5rK9R6Gk26V+SKHk2JlbJTLiWoLsxOX+8pqGaHnsPg6Y9KjmO4leU706VHwIedbUr7
R9KmfeeH6S45tHyqcQ84ix6gToBReKUGM0To5+nM5GxGzdFDKcauWDhBynSAcP5C4WA+sNZQDA65
spPYRLbDFnsMDL39sSY8o9HcNH4hSmpobq3MrChMuHHUBfvVi6UQPxHOwaPrMmMGC7mqB6kzl9VO
7W7qm3PKw8/Gv6AiRwUCMg58a/tH8Ogvu/zPWaP86PU/ks6oHcwIt97/sI2+eL92FkUbcobvfkF3
a/Ype34vWk2bNIh1DiHAdXXcQdjLM8kZj4oHVU+MPp87KgkS4D7dEZo6puotcWJs358X2gESXbEK
mQwuLXFy9zuHpwjoyzbCcfpVkDjF+PubHil1RCiqo0NF3M68y1OA9b6NslZiJDZtQoA4+r/3ie+K
UPZh2NKezcEakTgRTP3luYv/gVYpG5hNv4xs2ehJZGiZDDxBi96nDmBvNLow5kbEQGkFaFPKUaKS
/sWxd5gq9oYqSsMMqu+2enYBhPuc4wSr/HH2B2PMKmGuoBaafVtM2b1xTtbwrGiFEEXsllwLBP2A
Vi2LDfPpCtl+dJujYUFs4eQIwu9KrXIzTzUA/ZS5x+pmxCZppRwwOUVajn6FLHHtnM/TftP73sUb
PQTLqmG+bBqWlEEnqWGytsHkh4f6JlDBLZC3AYVF3zNHR7QgdWcUB5LZsc6fKPkzCwXrDrTFUX1v
y49jku1WDdwhBqMHvb+Ou4Wiemqb+yT1EyVC2drsZrpWmx9Qivv7cnitT6622jdz2hBioyPTbdlQ
ixQ9mp/K/Oxt3C5MCCfdcUWdedvKto8N/+gNI165KEoGilll1NHH0p112djOO15qSV4lcrIPc7VJ
ETReXFe0p4Q8e89OIXHRDzQUlrowslbfufkhIYWFnsjqiXsIEF8YWT6Z/awWV9rRizoClLlxEdqb
XqO/MmkJ7fusYYJoLuA3tsXdUSujUNlP4rN9RzUjgL4TUP738O4zjTFhrmQpmOiuib2p1/04cl5j
CMZE1WkrnZlXpXclZYt6eEQblP4/4ktxTiQeqNtby41oI+xZOSafT0iqMifuynZJNEIsYrCkj1T3
rb7ZLHL9ASrQDGt43cJw4s9Rs7+7Vak45mLWK1zfWIUmdtCYgCO/Tf2me/2Kwm5PF6iF6UPlUVeC
1HP60mpkLbeBFdOZrp2YuERnI6S9JqALnqR/StIslUn2V7+ZxLqic3yB1pydm6ILixuTFkPgkPVD
Sq4XmdvT0Sb2ursbgOILgSkNCEqVI5orLyWXq2jzURAV3sOYxzl18w/3ydgMZnsppc0SWy2kzOLP
/zvdWbrFWGJtd7YOb7Q3WteUYOA1mpzMRjUyYOFpAKPYblCz+WuSOWYoSk68QHq9FstLca+fWTB9
eNPGUWZAeJW3kV8diUb4py6lcVEnSEA8xmMxWUlLkZZoyeMM8Y7IVM8FgKAq4AKht6oaS/natIJE
gkBJJWEAYXd+M/DB8lCxZbQSx6XMUsQIFtSn235NzFctHkHpEUO5+eNO0wuomNGpH+ICGuKte813
8b+Bhw+1BkAtgmgscBvPq2oWf/2Fwu2+lKRtWzSPuL1Cjxa9kT1t6rQ/a5ZlBENhtgIRtn5toGui
OAdCW2HrUkgd/vlo0agetX9ENOLca6ByAUuqoaVuTbjwx9zoFmarWlBb3Oaa+WlFP5Nn+1QJ/VJ1
QFHB4guPrxuszjKICj9XlVYRiKOvsygNBKJn8e4KCjY0OSmudHMuKXvjEd2+diVdmwa0IipzViGL
hWJrj4OzM8EtbjOiPtGOJuPP+Wfs9hrd2iy5wD639tPD+NWO4UrdvvPImvF38WCTsVyPM6ndmWHf
2JHUsB+R1I/74ERtf/50ULms14R/idl/Rkn3zswxt0QDkQ6ZwwDwJynIdUe3lpycfwtFk3VqYCPQ
sT9K8kMD2I3V77FwQ+FWdirOzresHOvzQ3ltW9o52zLMFO9zdbeVz/H1gAR4vL1rtYIFNahYBixZ
UHRmseoXfiKJt4TkCWXKtLgjhn7sE1q6+z3WIi1u6ZKw9iwZFSTq6M8avS+djlVIviBh/O1AdMG+
DyxKQfiaDLDetXPHv02vyvTYdCCRiBYxr11jfVvDF6AY792Mh45RJx9iJYGSjKFxxCsEHp0UltzR
mERj7/jjElKB431e4h0Zg49uueQG8NNf3lNvCnRl0E6BjvtIGNX7vab39NlTq8AOS6337/CG9e1+
sW69qvpOsErUdoLp0wWWStqfiy1Q3xEP+bf9SB0WLEHpvssgVgLP+d2bc42/GoFQ/viphxRM8Zwx
dEDhyYx6wCS+TGGapbsIjyGVVLGmqtdA/k2PdMcuJhLPYxBFj9PyI72BlKeBew4rTsETmn0vYJgp
NqL4VXLcLrlQjbzpntng4ZGkbXaIYvxzfg5URcahys7WQLZMbDXZXlmancLr/Xl3Wk/37fr83Jeg
jYlqMtBpyu1B6dLUGBbK2EyZEoyvAYQSGH4bVvOc0INwvRRUWHfq1/qQjscO8BeIETOJKYYzom22
Ji8pldQqxwPaGWfTLZIiX27dcLnIav6ioEjfxGa2dWt7mqk5M0C4pwEPjYkeBx+VH8aFCHBOJ4q5
/E+2f8KOTGPeShAA+SeRDgzZUXhuwOx4softWF1C8cBjTlBhP9pWxZXSnuV5b693/AzO+18gLJmW
r6S2MIfIPPMxeoqOfJemEuNtGy6HCrr48OUyrnjzEi0wRK3fm0qXw7RGvBHu3nCeai5K0A1miY6j
r+eeKiD/q2A2ENgNVi4Dzq6hUfoK+/luW2nWrr5jucz8DtEzQ4qxeilDDx8rDSu7/RZtoZEUkgh2
49BLWtDagbphSnfQl4HRsvTTfQE0WuTXhyL3tY5B9gQFtU4nQ6oHSF7nCrh0KQtFXudvUBjOEO2e
aEnOpjGRasvQ51KGTZ55i5Vz1mjZoLab4qFIEFafAJdKGJEoDaDU4Ee8pI5Pvy+ym9+Fpb62etnW
isl/gqestJPqBterlbnxwzgZxKFqFVJWmUwAtcDD7oJeDq5N7X+lrbvVJD9Q3gCjg4CGwz1DwSDy
japvDCSUMtkdr/ttS1XXTe8fBvFpeROojGLKFhJ4FEXlyfVGW8C0JBeHhJNfmFxzuu0eDaU/k4Bv
79rX8nQc71lpXQEJtkEG14cu36h77qL/MZkiOYQQBACFLi7koCNz2FbhSdKIbV1yUA1jzFv1VA6x
pvv4UFKyybYiEqFNnIPoc4sdKEgFUhoY0GEU76g0FOydIZoWyYuoxZLfsPchzQ7ep1P+8zpBsxxf
fB5yyzH7m80lxWypeGCDoOgxi1nRrJVIRLUaBOJIpjd8BvuFG0BkeUqU8X6DA3YlVAQc6JbJQUWC
rcl+B07I0fwswK303mO41Z0YTOLEE9Ksv9OAnyb2CA7Mms+h+2jhFKyV4I14umcjtS+HFoDXT0Ct
BljrnlrzMsK8ksMPkVlzII3QAg0eEP3UtJn6Zc+xI7l2LbxjzXq1olrKGDZrRJ+0Kjtm2dwskilj
GThjmSqLitU+s9bNDkzh2RnNpxioZ+Qd2WJ1DIfROQq1z8Amcc9On6t/7wwjLrGQ2Cpw5Xhs3T8G
y8xTDwHkuKaiLWtqXL1H3DUUjJBKorVbQ8QGATLteB7Za2v7+gvQPfRs/kBf19BJvGmq+reI55Wu
3QZSpucJ+ZVhoNT17xHXwO3f7iouojQoxU8FH5mQAi9BpPh4rV6WI+TDTmH/Gkn2NQ0XsOkkIiky
sI1miOC7ZoSjY9TH4RzzP8nBXJj9flJ/jQhNg+O3IE9bdrctnYB5LTpJikvV1vnYOUl5D3v8IjzY
sRgN1dcGLD5hycgIQSj/lB5c0YsgOcT4LRkTxKv4c/xHMgcNh3RKE3TU2IVE2xOdtdXXqEAHDsw0
rZ/0vZPZmvOEqYlW56D1dpVhlZ3bdd88ZycHflm5QKyYEgmDQkZEB1p1uUMNcfsCPAeGgOTOwhjP
Szw700JpMreDl9Et3ZjKB2/HAPUJmapVV0iARd4RbPnHPdUhoCFfyEQzzOUiHHP+fL3Ovr183tHo
zQRrlXJ0lpeB/VEX2icfgtkgH06dyHr46x1Z2z/s/fa5ITV235GzL6tZ8UqEpZ5IiK5COwROIuXb
TDqPJJcesYpcPenxR3I7VzJw5U/VnoWRXyfDPeahMgc9RdORfqBJPZwvtn+W8TC6XYt/VC5HX54b
zc10GD1wXHlId7WKCz14kbsYIa9KVanWhk0ssiakXERIcIzaNKbgfbC+zH/HeoCWmfnLAFguaU8c
WVbn15WuSnsLNF4FYnDS9snltAIZ6XYBfmvnoq8bORD9xLHjWebg1eIlyXgaPTaLyj6+6jjewqPI
Oo8izbrn/dvUVTWMARraXGetzsU4B9baOGrWQPviBliGlkvIbCI0YlqnL6fIbIuzHxhBW2Dz5PaA
AKCxGTi/iyuNXRUbDCC0vWRABOBiHm7n0tAMDfQ1hLLmAC//qmLFi6/QRQ+TEPATkGdDJw2zKJpe
Gjf5trNQX6MzAoiQSC7IeHQAQdd1cnYN+0JU/A4pISyeY+lFd4xkdLjw3wGCc+//jePrn5DUZuKB
8WUHbJsAGsai4efZsbajP0KqEL2D+lw6IZu/LSex0YsV72tR4taEpx2AVGGUVwUp/i2bKKDHrTpq
gyNaAZJL+VuIRxsNc4V0LpifY1aJNS7YOP70VRImGx0yqud/nQ9VyfySP8UWGE2KGyCK9CAEkFFk
kNGcIMyRgYR8aU3cLmope0quLMp1LuYLI4j0EmwnHIbEgSF2Vwt9ra+l7NXuhNGnUWm+FSB0IyzK
nFB0E6tTQZ3ecBX/yN0iIWwUwu2fiT21xtV/XUhbD0RxoP+C0cS6hmnsvzUgYxAraRj6tLRYPMYi
OwnWT1PCynKrcXw4Szxps69Dlo77rNSaObA/iEELeOJTNd8bHYmBESmvaxJWiMikt3q4c4oZQVqq
vZK2bT77lu/c2qjMuroVpQlr5nTvHnUyKaVYanHuuv378H6wTb9yftYhI2sPIWnctZ4BzZC6DTd3
H76mKLIQOYmL3J0utk4fbcD3aijI4YLvqy3aRN8X8HT1gLlAAEG41+vbmrdwzYyrR+Q6l42/hVS3
N3Nmzjsh120kZCnSPsxIfn31kSw3+juLQX0VG/A+Cc3khd4BlFl7o1rZopsbCS8I7hBsJmzgyvR9
FZs1vHc97iTPveDApD8twTEtKYliHG1yMTGa1C963Qj9DF5sa3/TpkmCIqgbCxf6/KvK0YwSNPWR
pQdv/GmiXI+KqNB05Q3IWNNYoDDdSzv+SjN2HHiqvwrGEN3TfWi6mv+1wKPdu+o20loiSdr4Tb0i
bJ9tQ0bYa1aOZGh7TKwAFIG3513Zj7Ob/76wgOSOizMBxg+FWJKGH3WhKhawFsI0Zpp4HUebG8hb
DVO3ZzVr7Ehp7cOcaZrfHZ1aAicbtKSs/Kxcv7NqNKfxtJVUdHnUzdqcDybxyjbcjWIFDEx2pttj
m+IU72jCo0UhPjjC/OexBItGlWV4HqyzHeBL3Ag3i98mrqQqc9X3aBMesd2Tzj14EVLSegwcQJ+p
NiLMDDuVK6oYOZMCYvIUxFSPHDzPoGfEk+IdQo2x9im/e5wIJJrWj6Zx9dRkOWbamMobubngwbtb
/uAus6hHQgoOgYUkSmtqdSnp9EflavnTQMkozI9dZF2cD92UzTdChhIKtQvaR/W/YbW3ACxAix8P
SXXPTRMssHztxS3MnIj1RukeOu7n7bNnAbQQ5i5G/kpDp54PFveWXlaKod0sV054ynlPtqkHMHBu
CkOeeJ6MuH9P9pVZUPFa6bsm+7ckeI4RM7ytVbM4VpxqjORc5K+nCQ1dTMxkh0pcKmnaf5bEuOWF
KiJytDCPrRBpUT60O5dd+u+9bj+g7mXSigIgzz+ZbbWThyRiteXlXsVBInJFBNCScqQwL88glBdH
1xEnusV9/kiwAQE5dUfTSAXuNKotUBh0klbwuiIZuYQrwnLFRMp862rgQC3JJ2jcGy8O8TEx1Qd+
71fWAsNS04VlTXDTCFnuw4cRqIgF/Pw5n3KbvwxxnQonpb5e0Mo03JF74pbBgDT5kjVqEqWll5U4
8sNcMRSHyDq9cz95Zd+4ETS93fZUIuTFSiaQEKJ4OUbJTXaYYUK2hXWP1snS+yOWoeS53WtxJ3D0
iotSMR8jRto8DYBSJpiYl/7lN0pKTtzT4Gfws3+xneGLYuP0ibiqPTot3jmpNBbzK02vJevAVsQH
vH9Cf0qCz9oR87e+cgcm2uVneG0TQHTF93eqqJ6jVNU2Hfq/XZvkhXDzXucX1dEvMt/Gq1ofC/7O
nkyq87NJl3YmXBWV+JxfMNCwKJrMFbv7CF+k1e0Lmh6Nn/vY1Ry657+700LKK99xOh9b1BpVKl+H
6I59ISWImXE8s3uzxRcdSQCO0DoUJ9IUFaMpwIpMNBr8LSj234ku8Cj3Y7dZuyA1J0nQipi397mV
qtmvFxDjtW4RQH5CYzEQTk2mE4Q3VXxj5r5a8veTyD3AzWWy3uJDq6bcIJWqHRgEY86JqZWA2Ar+
coNjStuR+QTt9Hsd+/VVLBns4HDbhaAGiZM8cvwZIzxgVdcE8URq5p/6qkUGVvWD14MXbbsxP2Nl
GllFvN6FcuvfW7NQy29mBI65sqJEi+9J78qrBCQTijD+N0SwON+/adtk2i/kYGR236PpO7IKkhn1
tGpnCnEobEiW+Vh1QW2DgGJCnLgy54Lr3q5S9yLh9jTpa19zKPhxKYL6GUuOHyFP5+GRPrs5C5Kq
84t8YSQAPFfgdCh4L/r1qJib4XyM48c=
`pragma protect end_protected
