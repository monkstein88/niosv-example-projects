// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qZcwDTd1ljAnrrhFj4Cxw4jGtPWHNR91m5DKnDMuBgP2ovog29/e+lrFGmBqnS/922ZTUS7dWQYR
ZVlfJ/xMPhg9obb9JKQCeDEI+fg5rzvU4ta4NaQRMQXHRxLjeNCCqWZP/N0f8Q0xkU3tG5XQu/1g
6iMyKc7xqAFZHICTKRNZmwezCs/WajdoC8nNgrkVzbm1JA1xHnoZBvVljs1WykYEMafhvnqz5Zh3
ZqbjkJJVf2T5hsx+xk6ESGL+mGUCntBxoKsGFw9q02WMt0NmbsBTiDfZoUXdmvHxSPzWxQuICaam
MWmYj2DGCZet0Iic70iBpb0jHZ75q3yyx+dzHA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 15376)
KKb9JH4xhUcbmQl9QKp3XgxOdVSmINQEkvXDMvv2e9ITPrPR6Ip2VdwfYwV7wvVPl2vtlIcfOSV2
y9QLDaIKTZc6cuY5+MtZ2dNojQE/CKa3f0BtBqwR0pz0eHWYM8SCVPSrViTxSL8YiyNeCiDvyNtZ
w7PSoO7AQL1iX7C1JxY3MHpCcXrvmvFbl9vl0kt1tNzrkZ67PoyCrQeTmKtBZr5K/9YB04L9YsQ/
1Q6f31GgxgOfW2oxKVj+znm7ZFnl+jHM+wKK2SzC11Ia4XC759FMrF4WMKicT5dt2Oa9zUakxGu5
/teMeb24m4QesRJ8rpR8mfwIc+UNwONVys9DJPlQVMnBa3us8xtago8P4OrvAkmSYq3mUzlO1Zk8
ssOup8jn9yde5WXvAthDWHqD/o7LVsEOgTD4x8RZzD2gZD7tL+Jv0XevfYexd5dxqKks4Bceqatd
76h3JEFPh/XthlNJVrIl82en9bnUONXCj5zXI09Xzpt4BnDwpARgj2xec6ZDwNl6kceimGIgdnrX
oC3D5en0DSfGGCGLc+Dr0/Ibi2FfwuXwoKBcKK/JAcvWZzqx78ZH0xNXf5GuLy2x1kbUa/r30ELZ
DgpbCDfYpygW2/q7o4dhhCjx5d2h38fCpAijWi9Hp7jcYa5fqmfp0pLUf2cjuFzMjJVeAUy9GLWD
IKTsFsy8E4KwljZGGobDYTQjaV8ZKrCotvHUsKJE9sbwXLEXLW2v1vvmGFMZDiDIDOdrZZd6r7I7
JVTuNHh8FZGg1HxSLKRyLgWWiEqePUOOEpdNOn9jfFurx0YZ6h6RlJBAWi6f6u3QSN6YwPI5RYsZ
jXhaPpwSZOoqrVzZBJwyibAVnUThLX71PHRkpNbGlVnSy2FAdW6HCsNoOdhb/6kdc7Wy7k3rWlPk
h6g7W81+WwFYwRONArQszLXpkPcoi211I9bNRPsTBmOBFpYviT4GaGrLA4VkS7rriKNKpHYk8Io6
ML2LVkGi8I3pSwJI1RT51lXqLYRvlIpUNx0338AJidArvfchlSzUTgVch7+M5JqziOf7QXx7BRlC
mXPdGTZt5GTBtB1puYjHZc8K+yrDiAYhDfkjTDpJKdMYceCF3p5aQo2FMlTjQUxUrVZs8J2TLSE9
P0Be2zNs2i+Y/TaheEKermKLNQleJONvvYMb1ISDGZnmvVQjmtvDwCwai9Ug/HbImPmOn7r/FvQJ
3vVGLWFnn0iPoRrLA2DQkzC8Xl3gLB1P1mYmfGG8qF4FXTsz2x0LRyWgFNX+xfydIZ+bInZX7RHd
3qKZn7l717U5B6GOrqCRbV1yEtMEysUsQquMOsAeZTpqIf+qNRnl9dfWyQAJu4wwGdFKfzqLb7hv
lAUdI8ru8hkBOFOTu4gf7yRKmaHqSoKpP1mkVdY75ypz+v5Pe1Vz9TuJyO50Ct3eyJeZblvF3mu3
ynlMSdr3S1HXJ/TlAHVcGLxV9/z2bOYiYoNR98a07BKFFgXqvUPPBlqHWVl17kmtCX29vfjmHDE/
hGE+vGchVpr2cA17/9gAfk8Ay1wsNF2bE3qgxMyRwcY+uClsfWpUnXcYhJ0I6kw089Nx5Q4aWdy0
BndhKvC6yMqEZU/xC+ZXBin14ItrkL5QG11EFMSw98mpOe3B2IsjJThEdHKBvKCBr6WZf5MV/Im1
gJAFKXEDQYsLaphV/O+qfkHx2qaqE3Oi4fTtRlid3PovyG0Dc4Vg7kD26IqQ4Od3o8g+CfTI0OhT
aZvD8WEfn8/Nx481sKhmM2VuLecepc5r6geYKmEePQJcXl3OtOc+l+MIVM3uGODPxClGBhlv+LHV
LeXXfnX1ramxrjHCRmMX1/YdoVYdcDkeQBxDRygq3yYVANOZb1JWQi5J8F89ub/LOYzIYwUS5/Cm
KHDnnWwvhMQtXVVcW66nK2tYJB1mYxbjdbwaH2mcb1UlRWAgZXig9UcTSU/jDODJyRhOJy1wvpBk
vKnXhNQjBM9PyAiOHDpK7lxxaA5YyiMRmxLRBFWAkvXgLmrvtdgr1j263DXET/dg305KUstTXUjK
5R/86m6wYNnVqn7vEuPaOEiCPqL+/kCXfOc7XPMU2po6ppUdgX+UYU45nbiiiCdKu4GgL8m2FumF
YEfL7i7isG60PD7Cjfi8xnnSnTeMRoluSOTIUQVeJdUPTZt0h7J8fxit0Kas4Gbz4uQzqj7OiIRK
YM6qiKcCIgKLp6HEqBmD3jlcqMtK4ErgUp4S+eeFJXYhT0W3iLt52pQ/JylYqZSYbfUbRnXKjsCN
Zb+6QRyzj1dFMLRnWmwWIW6TGazbaIzp+aAL5GAsDHNdgWmAle8Y9vm78gr0K4TMCIUckbg83fBI
Kf9YzJusslO5EjfhJu0Rsj90viVDSl7EgxrG5BKtrvJOTOTISjLZqnGWZuD4+D3Bv1EAnV+qAmKu
dC96eSHskPDpKU6VyRN3tzk1KonLWhhcE3QnDJJJ4ATDE/29bP20axrbWkB8hkeVMr822brkNqsN
zS21u/c3A4TN+SWvTE6JAFEVt4wMCkhz5mBax1goLLwHN4AsO0Q0CUzldgIGz4hfPXhTSY16USYI
yrvIXK/fxMt9sZNjFKFiEsC+ZyWTxl1VgzKENAdvMQ5dP9EcGEiGJo6wPf8Xb99KO0EiIXc6nuPW
AL7YxznbclfBxhdXFNoIs/paQ2FoJ3T5BgbKs4Za3fdd/2njZ7JnFonSC+4aOUiPuEzOZBNSY7u9
+4gTwLr36EcrY6JFiqu4y+RyHfUdIcSxJc1RnD8ldpvV+ywz0qWYEp7w0BqN6fkxRyQ2IQ4j9fUa
njMEOkpO4YMR2fKTA/ZFD5CZXrM2h2dJJ+cljqGNWly1zi7+NIrVCODX8WIhpwC5HB4Ik0ICII7I
t3yr6h+w6vcra816aDvz5+5swGL771GDUBKzQl9fTrtjhQhokzX5Vy/RwyJfeARnZlYRli+npJt/
6H22lP28tMDgSkSZVy3P6r+Q7hkVzmvd/KaELBAZ6EKIacDoekEydSXKzwrXyFjjvxcCmttJHVNI
NlaE2uLgdGRMPitWyfo4GrTwVPrLoHS9gvqDyOehfvY8YoLArDSmAyWXw5xDWYdcm8Q2ZLhOGM4G
a+Y5jEwu0tb5UCBhK7Kx6WBKYTtyAjm7ujMBlZh0SXAR/4M8xS+EPq2BP7inyIgQVCOy6jVh23jk
WImlH44zjIKsdtsii3UCIKlFykYWoAvk8Jh/vQ80AGJQA8eHuNexVTO+Y0++FnLPTbFCg9X2TOwI
xIZNt2l4STAwnsRoqzfm1G2zmQQF2qeQqXb7BK+zW2ot/RqHx2AaYBG61y9DP5ayo98R5jlc4TFJ
XTU8842DM1xKKVLMmAgK+2/wXi2Z/yPM2Nf6UMCQQkHSYaGfUYLpzqOX1CsbBosvdHh+CK+9O3Ui
CWRoiPwoC6SWDhI4OnLwe1xJ3/tqsbycGeF4AgY78WSHmjTPwzpNQR74+RQklkmY5EIPlJBuAFUz
wAPljVnnelFT9LBUgiq19ClUa0RcxJ5wY0D+dgE0vZuuZGV+N3e+hk25qsZspXyzdOtCM6vyWzmb
OKS7sMkV2KYJna59p9sfx5IH7zGpEbFqS7S5OF5XBNWcgxFrOwxvZ9CBo7buVgtiBEzyJ6uu0SkB
dWaYWbsTT60gotR37mU6+mqeCOms9J4yV8+wF/3NVty0Jfspvf6K+7I0RpQNTdPMMn8rX6m1gqWw
4OLacdpp3qC+HLBYaBRwSXCCMiuQORcMq3lO7+IQvw4I2bBeZbDq23pSSBlK385JkwNGtRgqv1VO
ZnZ59u4gzn94xRXy1nNo5HMvW3yLvKv6+HFaI3Js8ZpQ6xhyom8JaYCAJnuRvsbW086cehhhEMkK
/ehjp3pDWCieR7AUA01/vedcyhYBF+sJx0pYT3DorvXBv71CP1O1SST7sMzQW0GlZNzuWq6jEcj8
qD/BO2qXFcFBwzliy4ltSu2jI6QCdzS1/A6aEGTjoQNIcPHm/IQ7PYnDR0qCw27eYheIuvm/TISK
S7dyR4N+ByO57Yhpaliv1NohWWp2m6gNeerTTTH5iOGy1WrqNUyNnQ9XBHtMHp8PCTVZkA6z7jjv
stTUwxDmNVbYsxnBOckZVsDuaqoRjspU69gydUB/fz34g8ki5DFXHhJdGj4zHkBWZJXXCztQENOF
CTZMpbkV+rxE48hVi3ckI14AO5cCTHqlro7JY7SGNLsnpBSFk4PLHv4QlTt0rj69a7WZe6Xm3rgM
rTaA1/UkZw8IjfbhmoGQcrk5VuwZJgXCdT2L+kjq4KEWQpVf+/8mSsgbSXpFXHE2q17EovmT8NE1
IOn8d72RdTf3n155EuVbtKJPg00d+sLF1Xwphm+CFaEKEywIhAJqTc2tthKthW6Ln2+wF3z1ZHMv
ATHFN9axNdfsr/GquyDbapIO6StfPq9Q9ssCqPtFgolXS1h0n1Ln0uwq7b7OyQP403COacdtFZ5J
6iqNTNKdH3fruk/oQJpNNW7CWZAarbAhev304pMP/cEDGByj1CdafnMwax1Iueh1FZMvCzRdSaQP
EJGOD2zuLtJYynAw0rg8cCUeQvHa/vupXnP7epVtttMoi1xmbmsFYuKuKyfauDw9dV19PCtBrjF6
po42xMEVKHm9IqKhMgYhq3RpasMNnmceo+Tqref7/dCM6asWnQ1YuxuQ9k9vAYnEEj+3YSdgliAH
W+txW+KvorpgVVjytHhtXAOHWKZUibSANSP0MtQzbkBS8DliF7Rkvl6JUFUacpwSUfreamxQP1Y0
CrUhmcOPNbEVcBCnT6JfPUc3i0l53vmwb2yuDeXeSgXMFL8U250WXsmX3aFjJGsJIVvafSmD44H8
LwSZb+lEF1RI04eH7H2AOehIfxz/a3b6j+XOkHiqXqcCe27gUb4br5ZVFkYgZ/d2tpk/WzhcGEEv
7BDgQovj5c8hEg72tLrcgCSlMXsq6Pnk1D3Fkq9HgEC+WPQoWewZwjyh+I6wDnECUa97YuCxeGgS
oNLuUhLYwiMMN8OBaONqG5QPZ+D1/piCbqUHaryVSdiZhnSLnM2DRM9qxobnCIhnyt9Nb/GdcpJg
q23NQ2/c5MfjXoSLsgy2u9kZ6OThJo8jWA0wAjPIGxpkRA0mEkxvhk8OZI7pLXjgP0MCkE2iq6cl
c6/Ciy40rAUtFw2dRQAQNa/n6HqavBrlJNc1vXlpE3OBOEh4G/lB5wIXxPyIxlZPnyrBCjWH2L3k
ycsRY9leAsKlPCtFsxl5nB0gpyO8Fs0YyTczfcdtfjeWEICMpyOj3oVBUzQFG2me6qaVE5OMLgXN
uh3dVT9O789qTPP80Sbaw+u4HuSUBgrcuBmcGlMwTzdx4G8D8Um8gcj0CSdRGv6pGQ4YTeJIM0fx
18uOR3zjPQ4HmcTpnSsm1jAVegWyfU5g771sP82QdBceFOxtjA3KFpxtgqHLxEWLMY1X5eloEr4Y
DXocdnaleg3bkm30Re3xBVrv0OIp3exHptLsnsFPBQg11l42ZaU4SyMP9vUEqIRp8ay42C1EkWV4
bg1y8vOWxwM7cI+UgDtUj8BzAbeNNHkblj812gSKo0sJTeXAYz0uvyiyzD7FYkcU3QG1Se8nRjyb
1dKjkyevJ8C0WYNCDbnCK1DSriOQjJSckcED9Xb8Uel7B/K6+iV4KWz4lj97x5tavs86BLwM4oqi
5vJykNdA7SBAJuobg2ARu71rJl4/e/1PjYORNa/H8MH7l/oYOECEDYad3Ni4tn726irrYkdqp8cH
d6ZqITfcHL3CGtK+8UnshOoeDAbrfSICA5NlNGExQadQCXoPXYXIPKzrqmTPD2fu4HgrE4BtqNT+
5G9VgqRv9CJ7ugF9d1KCh6aEHmNrfW3d0RLVjCnAQefLgegz+TwV4Ss/qiCs/xZsT7tg649vQt4e
gZwnpodMwIaIDKRNtUiUxAiLszIYGNrjVWxPoQsf8eyB7Pzz+gnR0Heqft9UIco2VLUzUR0lDgoz
Qs8i9kcglKL5d1ectJme5SStC+JpTxZXqztluep+RCdkBuLrwg86xzQKLP/9UdICQY57te7c3L/h
CNfejL6pWxvM28T0wniZWnj1hpR0EE89MPN02ZNIjFuJ6hAPW9Go09wAfFXYs5Co2dCkHtbXHPsE
gO4uN5idH6fb6Atmyz91ZSKJEPdTHVlyROHxeV6iGxnUNATlhRs2B5xwWB+rMju++I6Tyx2PyzL0
Z85S4Hy/Oympa50MgocMMP92rzi7EEa+VUk9IyooWojr6ehFOaCmgQGcgkisr5JUjlcJC+QqZlqp
VgH9BzZbkGS24vN015w/b5P01xAsWusLgYorQarbPQ/EXYjrSSHNT+bFsTHVb/4OFKOSiKDnUurg
SBU5QnenOa7Rczjf+IaK40npBxImCdvX6YEw9VSccSZui/Vm5WV5pgRe7sB7cNFigqJsL6xJ4Y3A
uC3Iyu+oclTs/1pbQKiCjcItrY/kbmkik5g9G97S+gAYxWk5XMkwVNZ1FmgsY3lUGYwrx7rM5ui/
zgMs9hk0mGx0a28nYIgUSrfBffDdtJPnet/zhlHQ15CEPVp1B8OIOcwgoNg9kkzB0JbUug3HqZdk
WLwanX3rRBsZFFz9uia4ZlLCtDJUl107QsvP6fp90feHIZjQwVkD1xYppMAzEAXjesJ4sSu5QYOn
OGUJWUbwLaOdIS42dJ4Jk3v0yPFr/l6WLRcGHiYOdmZlmkJZxx9EMAt3sm1+ozQXIIwE0eTBSHR5
6rRrJNSXUAOFv9BfGh0hTWW7UaBQ4l+UbCb/vrLQQjN79PRQ4qnIj4ufahaQ/a+NCGt/6b05EtUu
tlfEOGB9T/kzAVC4TaHr3Rq8Own372+y2YbhPlH6qNGkj2XFMNbPfcmS28IHeKqaHTyI8WJu5u61
9A+xeZiAGnVy7iSO6q0An136911OTpexprKDjLMD2zKMvN1Vf72m8WJAYeY7jklh1f4FGUSGzCsS
+otnvjuDmh8Mb6edazDkoKeDRyoMm+6Dpq8CTNlH0s0z6j5P91pJR2TxLUNlg5Gdmt42kF2CR+Ov
XHtZnR0jCc7VsgX37JAjv1jtk/ipV6YRKh7Sj0Rdo1csfopPcOdj4VKTctbhwtjRi+/9M0upql53
dugY+s5ra1mJh/3csz2ytDGZiCZBB7PYy5RSvPYNjkMRyd32gNUsrr1YZ+YANhDkifON2urwoSwm
/8uA1SvOa1MH/vnEhbRMQvYXPzwmqKg08edcZAnDMEICBIzQAa2n00i4gPRuJ1diNeiOtdj0ElHG
TU6Z5JR5UfJ+Ocxr/YebvLxhIQacyKuY5YGrQJoCELfGF4m9LnjYwgbz3OvFLLUFCDrBz5GlGV2C
hU5/y2GR+cR/oR8h1pL9bux+SAxpsXTxmkYPX3RuR4gF36M2OexGbyfJsXlp2pSGxfZ6/Zme9Nyu
VIOH/raAxVCGoTwYC8319tcfanS9cEvztkgbYagsFaHgUCXrb2Xvj8w6dyvdw3pynbfWbzT8s/gg
UChHfpQFJhumSRHj9gr0RIK90eW0R3aPZ6JsbZKG7DJy+0pTj8z6/8EQpElErWnbvWEAWrLBihQx
4A7hZ4AU4OVqGLFZlgJPAZDC5F8XXhM5KBXOOhVi8UOhZlv29s7bWXXuNEM/LhUoN/Qr6QVMpb4M
+RFegA8Kecnu/n8dz5efqFGe/wfzpV8xeUEC+iTZpt3fFUm5gMbta6YCk2zw0o+SU2TX0sQrbvmo
HCtVGpG7LBj/eVKZ1p2/XDNlx1klSau/UYYvr4SDmYvFrba7bZJf5R7wDPwTnY7IGdNvHnw6ULvX
DUYiUugmWu9vDNMLrejtIkxw3n9VdlmdhYGUwGLwZK9zIwZXTTKSmnoCeUmQpUSfQx/exfQndRuH
W91iun9M/m5JJwzcrBnBenK9CQfWtBKJzW/s/d/PavFsANmQPtEoomj6HENR6R6ygIk3oqZ5ENAU
ijQ48mGZk8MMarvdbq/8rqr+vP2Tc6A4cBBJ84hmL6+3gjYeRieL1MUTnjMQg1R2qKBMs3TdY/JR
07iSbxW4Xj9bsbYvDLBfFhJUSZJd9rjbYA5p9HxwJWcI1UcN0urzwh/dnmGWLUsLULQNi+49tZK4
btnVpjt0j0apVoNAvF8tbwYNIm4XX6UHBEFtOYKSUslGGoXo9FMAjGpp3JOuO/vD2o8JH3EfFmHK
eJ4/SZaZW4ge2nFqUicOPUfdfxgr45ICC8hHGg73pY1ninB55lYkhNfsGhnUgbPlRkLAUC7A7U7x
ofJc8KvCPxAI/rUvevsGOWoTaOkCNHVyFBTg1xh405yTELiurVJNgNR6LtTjpKA8uWVF6pfTsdrg
jNhcH09REzXT+hwUYNdYgGj8+0ybp5SkJmG1wuIeVtbv5xA5BfpTZl6rWD4/HLQb/sw9NLwIaNNT
kxYjniYVmUmGHceg3FWwpRlI6ZfWSEB9QY4K41EhZ5jo4vnONzHhqxERQGEK+KcXYrDcJcjO2mMT
x4gNkFXeFhKdW68Xn4yFsoyAsCrB0HzZx+jDt42iQusEwoOdWcJkP1tANttCPV+gffqi5uAxvRcl
1RxMK3yUUipUMtmDa1bZYdYDtzXO+EYC46r8k+qRPbgX8LgH5pUmxbOZVvL2UO9YOnGKE4eQa6e9
pPXbZq2RyMY0rmGiJ/L+QdQGGfi9Beq+ZcPveDTSCOL4BZELc2dLruLTmbMvqqYR3ao5JrMPefB0
0c7FcgNfqlXiAnCBfFXzngbgZVHeG5yX6zkHnv9/3ETaQheMuAFxxxRQwUuxwoKIWj1w6vZVD4QA
efrj/jPWVV+cEXWbJaiX54E3JUYK1Jdmzx+X/ASANQsZwPcLB3gKL5atJTsYKATHOdaUrJDnllG3
OjNzsgtf2/AK+XOu6rOD5Oj3uLaPJ0dchRDsaXKguKLXTMJ2oi57VcW2HNdj/BMAb6+az2VNVOPE
La4xC6lu2Rn23UWVmmtEafq7iihIEWd9TBg0R+oUlvqD8e/fA60ChDVOyt5wwo12c9qrNHy77ini
vZ6J7LaDr5xHkbO0pJxKgFPZNz8OHyYATbpuZohy+asdu6GVCHdFCiWUBEKjQpdROYma0x05su+V
xtL6evLwZu99x1he7t41vONMy9Or1OU5GZKecxrDLwP/AvHtPLkmCL9L8W2pAbR0hRtx6FK/V3u4
AfWawipLPwkDvPI1NYbBwY8fOrk7ZipF8PXq5gwRXXMLfhnNGRymqSZ1Hmo/cr5IkMeOaazIMR+H
tvFcyxn1hOj/PvmX7w0pewMaPp4a5HW4zqMHw5uG+Tb0Uby9Z7c2NcO8ZI649DSWQW1e56jlorsf
oXVbYGbjpGsUgCebonDy3vFLwIj+IoUOnZtnr2GPNpK52Q4+9hOtCXPzPHZhwmabxYbGuoMAua/J
aGSulOxakZpFCMUA1nxu/31arGZ4/Dv1KN92/ujNjever9ciNrZGqytGHuqKK/ppVevfky7byL0f
gxHLEDNA0W1c49/npij4Pwp8Y7t+cW6ZDgREjgixzLOvSWEE5WqZfBy8dcaG77Wn8nKeovjcdT6d
UvErSGL4cGmwhXU/vYcfkErRpjBhuEkrdh7ZE+paLO1LtRSTLZT574hs+MLeEy3IVux8kLt0GWS2
tDEFnuorwZuPqMMsa0zjMKdlI9tIxEDMNBw4lxn8P2QidBWCmMxjFrarnzmS/Py1sBnogIlsV3sN
OKHuU/PjmbmNIGtWtT9BFM50BGowR+EP9NKWE3SiIjlBgOYPANeE1XsK6RF9gGvWj1EEZp1sDRyR
2euT/GHBGPnQufb0Ni7XyUSGEqbPRSY2aZCYTtteR8BcPVqT7P87NaLgpcATlMkm5ACxgZ6EhMcn
dwwdW1+lplZsHLy08aCiTm60jBiuB/5gimneEg/uwrIiz6bPSxwYTkLI/3vMRReUU9SwJjDiqzxy
/v+6OzhWTY0H58IHfj8slNF7RRLjDfK1kmhVbxIPp2x0xRIaO1psCp7t/9DYkM7w/sLfLd8U7tJA
IL5a1LF7ZtPosnG1B/CkkNRbaRp/ApGZmT9UC5P/ifALE3PpnpIrf6kBBH0iHOiWmljk1dL5NpAz
al5e5DoxHar8sEj/pRM21zLJoDeaEeg2KehAyu2nNUaLDm2DepGjQX3UvJRdH8AiOjPk0uR3Mh19
+tmZ9FGqbBkPmNrZSvrgsqYkhmA0mZEiVqpstB8B2lbePqjAyHzECkkdtYEFCVdzR645+AJcMb2M
StUFevn1WS1LNk3v9iXqjUL3KqaP7WrDdY1n1705XXfY5Uh1xHJPHR8eVApUpuy2h2wD4qm0N+49
GdlEq+lIKk4X09GRsKnttdnYwxwpVJyPTaGHdSsnqkF6pcF+rsdONvORbXr6T8sjnqY3LHPmjgLL
2XuTtWS6GxoeR92IY9N87eM8UW/O/WbiNg7Rpb1tgg53taD8t806sfcfb9vIKTDGhoxGwEutf7gu
nrxsu3oWX9YEUld1dbCCsFSvQwKQAHFZXQcJ7FX2zEKDnY/fSPnre1VXAli/d2k1gF+HNxtQA2rI
WmkC6ejp2KxQgHgIIyU8i+1U3/pOScPlXMMKZIvFbKZGpkY4GIvK9gDQ7vyi8zGS+oj6PnnTt+7a
QvB2xSF+6EG+v5l8CfvrT2CLILwxrUWjPuEQSEPrV62HgqXOz5jbK6ro1UnVufbwOhw46EqvRpE9
/4MsCpKTOPLcJKVW+5tNN5EZynv1c/z9k/AhVqCI4LxuFvGjxf1Wf2qOYRUawQ+1iYWP9vgc/YNS
zf2rUBrIHGDZeSCci4ZqAilJ4YdC/6dusQ0rvSEsp5JBlbWm19X9Ylh/5l7DMBiPCJo++AYQVI93
+UEmeuCyvGzDMq0MeS5OQboKDvX7jbbr6hCgxsRb73ON2CvEw8bZHtv4RcAOwUx6HrkuvNcDhOOj
a8sYUPlApwQehUKJBFqQYkIxeZBLOnXSx3J39Vp7ldPIXefny1s52UG1GSuWkpfPirxBW144emXT
QW4p+GdJnO7EbSeMFxxJy1MZLZyIzYtTMVfIp06DviYXef6cjCIMiw9TMcG05o5lUGOI3MaVQ/p/
JFnKOjqtRfXKs13Jr9bCjWUPGGkEZ6iwGu0+wXDFdcm0Q2pTcAKBEqNU+UuVaNUal+krQq4FpTaB
Kq48/ywfTul30Y8k4fiknl3PTIK3jl22Ydxeih3JOM8TyDMdLxUHmk8wJN641YhRBOu8OGTKjzXE
9OvcERa2IE9U+kABHtL6/eCkcg0CdkzT2XBYyuRyBWITUu2fKJIO5/BzCslvfkAsFO7jMWjJUYrK
Edf6JGb+l8jgw9z7jhBO0/MU3blgcPsUkmOCkCZTwylUdXErmBXw5+LA3gnGPm/Bje4dAiAnspKl
Y00fzyOSpa1HlEv1OymFeFTd7Y8Lo3TjGg31tn+ZsfuVeCJGooIQCUkZLNS32GVaE2Sls4mAvc9N
7wTLkW02OVkWlU8TpJNrqStodVhy/AmxHNbiLKEB88rJVksjSOTXPiumetmOckx//pgHzth/fDPv
fUtuP0VLTPqTohEoI4tNVxlnQl7Gvd5NOMgIvywGeR6EWLXiKkTmFInfsnmpTR4QzErSNEWK1ME6
S4FKg/6GCgKvW/V2WSV9Ja1PvlFys4GBW604dNv1tyVPYtuHD0imq/E2oazmWr98LiG2+xhIDJ+A
Pi7QcAUDt2YO+TB9iOMdvuye4kRbWF6rLk4K/py5mrHaCdCuC3NrLO3Zgch4X7TfaCjV1DDgiBRn
FNip4wzkI/Fcf/kmEz2GfwFKtfkR7M2p24sCsXpzeP9coffDZQbZlz9s4n1tvXYUCTHyoJZYBpjq
r5D8IUJ68/yqvP9lHO2g122Pjgy9njr7BPZr3pSzrLRCMhhWSqKVbRVr+ht/wRr+URCYNK58CNUW
s1kLgR/78TIaKBBBBJz98XId9RRwZVn1AJcaahGm5UMRkpo/wLasj7B0degeFAb+unszrVsMBH8+
xSsz+d6eZBOGg4g3MMdUrQ2JkbhomYfsAt8RyWBJ1HGQRbEhvqcLS1ieAHs42C3kwun5nq00OGyK
+7j4OIEiKPFxEvb7hrW13xxs5nHt7fOCSd0TUdxYMx1KgDYw57EV9NvWafQQH3OuR1UdT0K8Ncv9
w2FGZjvhG6a5zBUJebYYhpzUfgESKoBQ4VLb8huD2Wj8tBWVxfjEk2WArJDeLfGUHsTBnYgWpcFz
8zdXcpPdqHzexsWLdBPIhTfRcqoDRcajKYj/inqqE8a6PLqYU5yJignYYc+VWCJPZa5DUAI0Hxd6
s1y+wbL4Hlpuk77ECLwIJQxODo6PdfYcdivFe30hfHBKLJ8hM/Ar2CIAr7+t+inH1mE7Zt/R7a3b
Poi+FyFDyK5r2CdwpbR53kfSEXwOtPfCDWl+zqtfsaBsadALtGQgvd0w4Nb777eh2L7nfhm95Hzd
pWzcylp4dUu4SLAsdmzHPp6OdYJOVpfBDvfOTqY8WvKQ6qVIgukJKVvR8X7xTqm3aXQuGkoN7mMb
wsdGbCeB1nizR8IOFckpDQfv1cJut9Ji9zOtm4ZyOk7E/kWxhY54RlPLZF/iRn7wWBuwdWK7URXW
tZF8K0QZMoi7FE3bErnWrWA0821QmoGB+CUtKc1xP9XVaphgO519sgX1pFVBymQ+Mx2Gv4wMxbd3
Jws1EED0Dxe7yurAXBVpn21xX7uwlR4986NwxQlFu9IZn8yYwVqQczAGl5cdB8h6k5hi1Igf26ki
mHTGk7DOwJd/IWYLwiLJ+0ItnEnUI1qpUEh+gxVucKOypWHEkG0n0/dcn40TIlT8eKc6cWojv4nt
LyGbCiwhbpUf3dDsj2UbfBc60aQUQoVvDAEf/Pr5tEQoAJBup5Jh+3f4DWHvUblK+gmuliFeIfOh
o/u3d3LifOYt95JZnxOikgGAomq6ERpxGgYl3/uNTFUSDJ6gKsgPzuCzFwJ7o/zkKpYRbAHgxfgT
FD/b4htObnE1ZMvaxP9sY99Un6wFbCpQv0/gmP00qOqcltzeMGYoV5IgLsgR7EIWQoQK56aZ33SM
sqVS4oj9n006DeTNtI4sX1VSrHoN2NIZfJ20MYg0FsUOpF6Pz7o/JhBzRjqR9WLAP+elz7gQTGbn
A9HVjl3ahX42sPblsn7gGDwDIx/nQNMbZPo2GpeKfCTNBApFp2iqr9obx+nhJknHzLL8KH2tO+ON
oFA8Hl17e7p8cQVGa14Xmr8l8TBOA12l0C6kVO4GWFISko1jbcUrCSyhUKL0i4Khma/9y+7AbT+m
vyspphFcftcjjJRzJ5jpn8IXJ1/bZ+sYAhlz0yxn6nUClhMh4kqpur3LMDQf/ChQ+OMmxUF0a6Mc
7ZyhS71lr2oMmB1uoMEBDFJepRtMQNIwh0a4buI/RW0xnu1EHCPi/QtsKmAe7ZEF18p/vvsg8K6S
KJ1NOSmFTdXAUqPBrfWh/p+x4z7L+cumapa63HRLoyWuCOYqrlQbiWnGqAZ6EB+/zDLOPjmZyQi8
yaumxSjPl7AQfvZQbvzyKoTC0Zp18thTr5OKfFOv9AEIYNVgGSx1rivrJQvC05df1shhOEECrOSH
dKvb6MbKTccvcJrEuICgL0QIF4OFaaQS5vjmGDMLoVav2OuK7cR46YeyBG31rG39LfZI6cULeZlU
dZT8o1hNKgoa2fiNwMt0Vmsn62f0QsqzQRsDcibX0jsM/RJhY5SVtxzfjW9NxifKb4SizAy4c0kI
edD5o1UDGoXSvD3dYvVT+gb92EYTvA55mxg33nfpsojYzP/+knEjPegO5wWiCu1cx+06KJif5kWs
MRgK4ZKBrCT1UAV2n+3E+n+AbsaxI49BC9O/9nxHUYXiUBJPOeVfZKoan53AitxPyi9JPw/BYecY
Vs3s/EsQAQgHx98Znx9j6d/BrcOW5OtckJFxl85JDdGU07E+qPH3lu1SKb1GXyihKsMZY654aZQh
ckZrhKTDOj88HxFp6bp2FIJQ1HgxyoSh2eOXYFXaEp/TcLmOSwntNQ8nd1wlLhs4cEdhsPcOqOoL
x6SyPIjvSpILi9AmjG5/3Qsrnv0Vdt1Cbu5KvaOAa49ob/dMV8CMCFiEZCHnul4bQoWV5xe6JUwO
QLAV1ZUIvUPzasSHsQ0w02q+GMen1Ibi3IAlNDNvLEXbML8AycMUHUgpyLalx0YJFe6AxkrTGUEi
XkIjGGU7UHnO2pd+ORi3mD3A2F7oM9kfHYGvSLjnLazLbGSqK6NNXLSDME17TT46eaLJRep1727p
RVNncHtPZvagrrL89hCx/zb4Lvkb3Ax2gzLXHsIU8IyNZ1hdl4hvEYOH57EWk/OFiv0megfCtxLa
ped/TvxBSAlZtL0J9iPB4tgXoIjFANUXkP3MRK0RJEiZChsFrEMLel0z5uf4QTYKKiFKgy0MLZVA
rg6W4kx4ZzS3zjQrFZLaD1OEyWuOqxF+cbt97OSJrCITowQc2vPGvSd5j/g5z5mxq+rmH+ZEOavz
rW8NTjeEupyD1NidY3AgnQGLX0AHZ72oZ247SJQk/Q8LHArQWeOeZL39b1ihD5UTeaD1ebbnK73o
ha603SjhjiDhCpvCTmJ5qLu1lWzTVj6Hz2rad9JjKSwJJTdfDoV1zQIO0Cf7z5/7qfrIXdyazL7G
iEQcS6/tVrMjXUq+7DUs+mUZc7zDXSKrNKE3aiC4bRsNmo2DNHeTDTCT8Fzfcu2wZBWcoLLb2vos
zpyTCZcE6Y/sPf1hgwGplQAQcn1p9Q08wXSsv+/VP2zSsIxVVPURTJdztF0GmfKZUfH4b78YMSjz
vewfPhXNh947QrJYMF7l8lOSwXcr8HNToRovAYlaN77gnbO8kUQn5n621EwC9b50kfXD6MVeFvih
tOWt9+cvx0KF7W3YZUz9GogEEZgOQ1yYT6WAp9Pcnr216yqq4gBDt+l0xoicif3Bv/rFXwqO8K5o
00y85APoh+oLwsBU515fz+FRMpDp8hs4ceEORgthi+QNWNKE9WRrjMfr8Asve/TttxFx+9eB+egT
C5jxS69PXN/wnSWuZ1sJyrjN0CFHjJa4Hj1x2oPdzRtuPco8vNrZByvtgEH9wkMHijuzCodQ4SIK
9dWxzi3buHNkGJbfUC0PUy6Bbgj/tVZmAWlkCErsAIpNFTak3dhKUcRQBJ/nadIbKelprlZo+tl3
yqACTao1w5UteVONQQn3pcLdaXwGyM3Ly7meRuoT8+Ny0tUhrYfsPPhOYLm1i0TGeuhVquuDNG36
PeRLD/QJFAd+/Db+GSujvy+OsyAaz7Yqql+soIfn/g9ZRwvKkXRk+gzJJ2e2BAlLSY0SqqGJzh5Z
dAHvksmNkmKqxTxmD8nySP5s+H7Wq664oJuqgOQ/ZMhR6YUjJqFN7a+pqsrm3AWftoJu8GbSMDvV
jY4hgmT0MSThpEz91jkc75QR7QoJnGcRlkwVkLH8WbbD6AqhjP8H1uvD2SQfaQUKNrk6EyLzg5gV
k57MPD3Lu6/eczX3uOsmfXgctSzoJncm47Ir5cY3nnYeTuIwcTjKjK2dCPEev7jTagm4fO5Idf7U
Ex1h/pG+aY/N8eEKuU9pt5Ewi7xdcUDbnQBY9xCueluJLqxVbi5LUN01PuAbBehMl3sOIbKKhOyI
LpXJa2lKMEiKcyCkZckh/pSz/TMdLGXVKO+mw6D43arJJhUYMpjHreiKipIbKLYd8xGQTQMbK7z2
APvi5K15dEWhlrhXuBSxgrecOOjLQ3yBX7RCzlRWXj4ky2L6/xHunAH1pJi2I7kcLyTP4WCuWl9H
oR3v83nuOuA3AdydwlPghVpcX0ZouBbAZ5C0soXxwYuPeYePEMgmbZsKrMRmAObKeZjBjk2EAsVz
P47QPt7kRODXSOkyZpfdj5z/MAVZ4ktiaXr1XU63AdRVB6/0u3jL+9SOvq9cGXCarZlQzirB0AJ2
AdQpR67zqUx74ttYpQ2Un3b4KuMZFwbmxVwYasQT5YGxIB2Y+SYARrDr8wEBjXJxx9+wjEzg13do
VGZ2potiFXQn+bvNUnzIeiK1Mfo0ltjhb/0xdT+uYMJcn0Wmn6xKX77fQ+kvb7Re/bhyevoZvUQq
ZKOwhBBHE0Lqg5Yauv3qfVCEPmjAQ2m9leRoI8XW08dsu7c+cMCFeULA4uAuwoCMAW17G6rOBoJ4
HvfasE+T+DVXJVw45rcR5dhD7EIC8Eo8oe1IohdH3lPgSYMZ1mx8FlVMVMhE1rT8NtO4NTDL47M1
yvldcJDyBQ952wppz9UdOB0DufCOoWldAe91dyzV3Npgg+tGNuXN0Bz05DyFLYxVAQmIIGmV4qXq
7AZApkIjK9OvWlig3BIDgVBvYWQ/BhLXVCdgUEwag/u09zw64gfynmxADxU1UfLLYOjRMqO110aW
DjT7Q2i1eW18t8eEms6N7H3fdfdGUvi/uj3RZd/StQYt8/ACyU5hdzoryRz4t0xB4yzkc5stOFRf
K9HOjyWlu00cbdIvzuVIZ+aDK8z08kaUI7R+yYzE4nAM/H9bILcXY+s1HgSXEquiUKz86t9LCmfC
rOr+jyTr8vw6nbG7MFnF19ERu4i2SuKap+oWAeCPRzfR0YA0Dx75+wVibwJXwrDPUuTVw6Y/9JBr
dQMaAVW2iVb5XWzO+jkzokphA9D74DDJGQJs9qMAN4ZZmY5GCNUXiYeyN31VRB37fffVVT46m6TT
P0lAzO6uQ0n5Bsvr52jnuObfEnmZQjzgny1tG5SZzbFcBCyOt0v5gaM5No8qibV/FRKfJ0CU0rX9
0G4r5i9HBWv0etcl0XPIF5iVYeDDfFKkHXbzZegHYhhFK3IrogrdR5kBL9nb09bKb+oSQFnas1NU
fvJvkD4NlX2VadHfCVqvxaf+U9dcyPO/s8rgOGmLW+00k5EjSkuVTiVmdjKNBr+B8MapAifhEdRi
ux3NAgTI8wT2nTGWkXZkUGqoLVwE+NmhxEzFqv9l3uGMrDD3ZYeUIDHDZN9cv46/6rAFFv/RSJM+
14tP5JnmbWbi/YzQWoLokKZeConKwYwnBlrhL9imCVkT6qlvA0BDkU78z+THtbK/tt5/MrysgRWh
Fnw70yUsaweDsO35Xzs/aSPt5NDJRG/jSB/tOjrA5FDqkT+GAwK+Lh0ogR47pXzAJdGA/wG4vDgk
+RXIkjfshMdeRps9eJbEFWMJZzjz5F0aJ2LSdqX2ekS4LVt6lNPVumoePnqaPkz8fJ1Cjkx1ih4Q
ZVe7rEF9DNyL9vChI1Mgq63AwfUAaqkiJL0VCQiERSAL6i0LIbjbVpg+/Jc9Ivf1M59JpGlmp6od
w9MN5Z91jwPC/tBBaGM7BWDIjEwWsoha2sK2avsOVftFJc2C2zDRfaumMhTt+V2nfZZJ94LgdMBF
5cFqMXDH9t3SVcxVqqCZfOGm1VEdO1wAfZcEa4qe9z+QHqQI27yjdOyP7MUzuC+9pSgCbtxXO8jl
DyBYl1D34xWvIQUOvbW/ViIhFrwxD1ai9zw95FZvIPz2G+5qYeEo/xufdgVaJuaaWhfuj5R+WE3L
TByT0dp4GYdfOOyWs64z26JU3r0Gm2cvdzHdl7ERHRxnao2rpferLMGTqlWok4i/U6It/IXtj9vu
xO2mSXWKvMhX0cyKlS123zalU5hHG2mN5QP9CJ6mBFmdYD52uV/zmZnLAEF0wKjc1/Qc1RZ8ORxG
auWLoJ0bb0NG66V7ZpKmG2tVXM2Lys2soLdza5wwe9I2Nnrk4NnaRF2r8bQ+NfOvFpWg9LvmnEok
taEls52ez0Jk2dgwuyqi4fB1GIEd+8Z8OUS/Hz3ShWeZkpYVEitno50PEjXN+RHAHI1u8up5l6iQ
Qqrw2PcaN/9Uj+tQ4rmMwrdEPRj4ZP3idgmVdYyfSaMey3p4HD+PrhfvBzz8L4vH6GTdW4Mw5JY9
8ALUQ1iz33HfaONOr9ICiHcAvfpN4WspAW2n8FzSGwvI7XfHttzsp4chhVJAUsMqaPafJpOV7Fmo
c6CUTVMNiO1yhWZW4CkGlmWGTprp2A4/V8B+iCVv+MQPe+MLc92XfIhPHdyUXLnqv4irw62pKqyC
ekUJNiJINYil4HsTyEWg49Clyu9brpDZc+1JxDWgIOJdAvZlPwgI5ICnNeMtN/0psvykopsikQcD
JM84srZ3urF5RHOLueIpTHs8OA2c/sdVr4zADab2aOh+XlK5U5kWEC3+AfWxxjAprlSlMbK73fKo
JE8mllhEAuecXr+H8H99bow7uGm1ehRINJkwA+pV27ZX2CSO0yEs48ifgkSYdD6A3rbYndIwQ1VP
9tLIYTQC6f8+jJa72fPQFiSM/PgDtiLsIKNauRLkL3k9ygrou8D/mJLY/eRpzkHOcQHCnIJfCpzu
XhuVgqOL4nEf5u2rIAYv7x5CfQvytjhNqlWwStz67efcainb2AeXXIK/4lQ1kk/aoQ0pszS1vnbg
+SCsFSm2iviXrezOkX0DctvdXSrswYRLsVOzg2xB8TZmT48bi4WVBXBTvm3PYER2NvqiO4ZmF66Y
08Tsbzw0UfdzOGQXFseFAhKGYDYwTlDiNuAVxhf4/yNjijZNQEwnkIW7DoIEgTYfO8Qqhao+O5b4
+XyTndob+rmOgI4QWO2qhRSH3p38MqhVJVpJxoW5YfJSfFkFMtRBRq9V/MSib95Jd5dqZGp0w3wF
Q8Qq3DFacu8x30W4mvSL7Hq45DjOjITR45i+hMc6Vhfdiw+xl5mG+iFspOvYDVQySbZYSXYmLOj1
gRSEKHFTR3wPs45lE2kGezZdKBCXvIywXaxXvUjkBv2ToTRwY5W6vQ3B9a5VcDGJCtvUzpo2Hni0
tK+AZ1F7+iZB8At1G3PAcSkxd/+Y9CeabBg2TfhAgPkb/HABKNBf0sWS0dir2yVfxfllqJ+kI9WA
5W4z0fzZm3cbcdWIn4lF35yy4lSXqMAuR8xiI3VH4PltyQh2UcdhFUclMJOSX8g2s91XgZyheBmW
janN7eA/fPiFh5gL7KL2wdYPNUbRiFPQfihRlhH0mbFLFf5Zw/YqISLgdYp0/QBpJfgKUIoWSC1i
LG4AiYs3RJWFFIKSu3e0T/2VD6FsrLjSSc2mwazpvWy30G7iwD4tQhNm86gJUnsKcWIZQEtHPwDd
XLDE7+Q/Ua6WOlmjGOx5SZrQPE6B3skGu34Iz7WcgfNBFT+K5EQ0hEHZJ98Ta8foPGCQYEJPchF0
+/L6s1SjaWuQ05JNNHiDONYZ0BMbpkofw7sTwBkdGQR23aBN7na8KDHIR7KXRc7eTJ5sghP3Ktqq
boRzetLkGV0lg68pyXhtbGHa1+ZTG5COOJbZAwhgtHtxg96knwCQRMJU81pFYCv740btojN2FDVq
4oUk9RuSRl38s/+gmfVIL0zLmOuv00Dnpo2skjo/bNw1cudynx82G2Z0P4irsd6EF2rSvzeBxOiQ
XrltaBtkbZ+n2GQPMDvIKA67wYn/xcyiGQ711CjjRpHTnM9MJEr1be6hobuhWk4JP4KhqjTIwrU5
Jq0s9um9t/46TOQv52c+kzz+bBI0xpECIcIfuVGxkDP0Ocp/eluPurFqTR5jWwmFQ92rhgTcTVEa
7wCBnZSfKz2p6XICHsZRpaA7Ol293+d/cs+P214pQwTGzhFEV2GTDU8jiMkSbmk4N5quq6sMNi4B
wYc2tQjDGepL5Kk2L+0lagXxXGkAoUhhM6FkyeZ/FUtMS7U+1WzleCnULx8HAElzNZQ+e7gXPSar
cRGDcPVrnaJd8DUk/46gmYT45/g6x3qQJgIXYA8HNSZ28T8WZ8ZIttEmfLk+lXMKt0yV21EBzk55
A3ADA4EepCsbDGTpse2ItjAW6xR3McqQ8FLMOhthuU3zXC9nF6f9RydZAjdBnbd9rNYd0ZHJB3CG
UM2X2c10HoaNrMklCJTz4tkxj8c9rZr8t6K32r/XSDKNeym/9EP01BT1V4dPU9i0Ugwl0AtJ8X26
U/PAN1Epmi18CW0QxkA9DyGGNrI4wXQEcLsTneEsxM5N+/tVA2dBZNhTp6MxCPu/Fbj1aRWrccJM
w/UHTCpysaeDn+GLHsa1Hl1/fTafbxW58+Vp/3L8j2qqRfnfe2zFoKTqKtWZ4fde6WmI9nKeXFge
BAvE42XL24hkO8RvRxkxfNStgK7uUiS788aOC7z8fJfjJ3MPR09T14yHAhEkFnIpDAZPLiPgK4EA
8R24/aX/EVmvJeyYD059sqy2A5OjOxrApBM92mC5LuezZsOyotILoh8bNqOeWYBKmbIwZyqY2xX0
KhZagKBVXsvvnulFzTUVQIun1P5ohUYp3en/auvYgTODj6+HUd2OQa42UOv8UFJhcQQhMtR9PKVo
6ZiifYPXfKY+fw1/WHgHubtraPYb1CTTXVuxHAL3QtZR6ZHKVocwhFlW0gYEfebobT0Cp1A7ru9m
tEhwFPSO5a81SN+4b1kjJUxhZqoJtGTu/HErnXTV2UXV4sOGVIPzCtbv1w==
`pragma protect end_protected
