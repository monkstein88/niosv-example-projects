��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a�����/�	v�+����@ɧ-3�����Iz�t�܀Le'H>	6"�U{��9�bEɤ6-�!�V��s� ���m�|����~μn���}�iԹ*VC�4���m7���-� �7�o�d�0w1 �⹺�)=k�:+5:� _M�e�$�"��O��0U̅�iZ��x�K�~̏*���;��R+X�="+$Y~�ml���n�H���K1,���0�ϔ���憲e'oN��D_lxY��^PZ�#�C�e��Au�֝��2ɤZ2���ܵ� �o���ǣߜM0ځr5r`D.ɩ�
e���
�Dc�����gC�8$����lc'�'@��A��Se��J�oY�\�?f�ᕭ�o0�\�O��H�$���m���M2�M��J��?�c��ˈA���~=ɮ�����D���B�p��;�e㹽yU4-����_8����p�R�C7�H��;v��F��5	��zMV�I�xB�cȀ�j��� l�{�I�e>;�IT�NF.v2���hb�]%fzy�0���#�%�GNאsXU�թ���*��j�5x
�P2V�?��9}��=�->���x�/#v��_�����J�N�(��x�USy��i7�4��J�ÞQb���u����V��i/��R�	J�,W��r����tx�E�r}ӣ��בrl��P=��������1+�&r�W]�#'`��5]h�?�G�i��:b�P�Ǎ�;�׈6����r�R�����
m;��V�j�w��^Q�Z1�d�p#��`�h� ����Ҹ"���'�1��o�}��d_��0�^$-9S������b�I'Ѿ(==� �����N^X39޻f�z�M߶�>m�84�G�d�|6� >��2'[�a[g� �oL�(Y�h/G���ܚ�ղy)a���l��� �d�,�f5�gFS4|�M8l> �����0<O`q�`�U�X�$.?@�S�xm���h*#���_��)��a��i��<g��Mە�����3xt�F�����ef̌�����:Pn�� EM�é�=����/�̣S1��$��<a��\u�!/�\����փ ���:�u���־��Q��2�sƴF�X�������)|=ZϠI�2É3�K�%3ń��q�؍o* t"it`�+��7��܌�G\{�ף�O���Y���L�*ſF?��i����L!��z{�Q6�BD&"m�"
��x4�n�_�������������T$�^��[S,��來d�[F�0zu��.Ņ�l}�71URVxo�]P��*fD٥��))KȅJR�9�F�C(q.$�D�����F�1���3�������ǱjЗV�&;�Ͽ�k�
�jk:�}Ip*39_�?b��Ľf��߱w�SHu��T(�������B׿B�
�I�%J%U��e|H���;L^��x��1��8�Gb��SV��G%�O�X�Ei�{1y�4��ݥ���1Ʌ�mA�g��=" /�ky�I��n�(-Ɵ��7���L�;��OK3G�c��M���o��-��)�����b�݄H��.&���f��5��~�ogwn��s
܆=�N=E����/�*5i;)��Q^����M�w�DW��IҒQ��n{7`�+�{f:��ڼNПez^Uyt�{ќ7Pǂ�	Yx�V�L�PLd��o�|W��HB�9�yL�f�Cy#��i���ϲ�Tq�xS]��X�v@e�icG��eL(w'�:r���u��#^��9��f��Yk�S?hr�hZkLm�3�����xS.��`�p��.KL�,��l
gmT�b��*�Pb|*��v|�-�/�w����%)��ծ@�d$@<O7�E�z�z;Ź�����Gw��N�����*��9�Z&h{��b���{blSq��f�dc�O���g��V������_1�r��Q1��18����7 D�ey9�p�bJ�[s�oԓlQLc��]k.���[��Έ`SY_�c}&e���V�*�DWgx��O������"A���W��)����(�n|���2�|ћk��o��Ǟ"�h��E
�̧�ah��y���q��,q�	'w����.�Ɏ�.,"��x�|W-' ���j^q&�����18����w@m�Y��O��h�0�'A>~2=?�q�tmy��ø��ʇ�'����X��ȹm�^��.ګ�j S]�l�q���]�P(��
���R�dS[Y*Z����H��ɀ�[�8?4����L��o�/%��4,��g DRc�'�;�z�	��7��{�Վ� F��
/�SL=�����޺�a�z��^�mb��@=�}��ŪA�;��9^y�ﺫ�5_��-}xΪ-���K���23�`��p-���[>��'�.�2Gwd�F0����).��hb�Eu��U[�Q"3t\|q�(�UP���,3M��y&'#"��yո3.���46��=]V�]�7*��Ҕ�k��]S3s}�92��� /�	�� �[0û��"a�j	5�6��]&d�M~EX�@��b_��'�i6��8*H��윯��k7G<N4�n�����*fy�Դe�^�����@�ʝ,�����Gg \��"��/��nԍ��R� �c����ECCT!�iQ�G�<!H�L�Qr������UtCw�2�?��Oi�P?��v�+M�OG�-q�꺒�*�G��N76�'�nKrf"��8�Ƥ�u��坈��j�?6�m^Vgq��
��
[����㝀2��аJ�}�HA���0}� v��&u�+u�HIT2K��B$�?tT��@{?�KV��J{��A�l0��D-E��# ��cyaOgH�<9#� 4K��������]~O�/���8W��?]\��w��Y��춹���H�<`�.�PV|�G)Y i���֯�V��`����|Q�k��|�9W���z�gX��vq\�����x�~z(k�{lƻ��D�-�9��z��;'Js9!�46��GW��6j�]��'���4s��ܡm��]Ql�I��������"�*lPG�d-�I�/B�e�5����	C������s!O�J�I�8;l�-N�2�x{��{�~�����:ĬGyK���ם��巂e	ӇOy�����%�w�(&��
L%~U����k}r�cF����ʙ�r'�?w��-b[		
�f�|ŭR�lhv��Ň!�ce��o^ʾs��4��L=��o�nS������Կ���mD��l8�E���lQjq H�c��o��37�N�׳ү� �����|>c��V�F�zf��⑺���w���K���f�ET���X"Jxm8�tRm��]�υ����ֹ���3O�a7�٦i��]��Щ�����h��R<����P���s�@g�K��C�w	�-����B�V}5!���$Vbq�o�d����+,Q�x�]na݀7g�o���>PUK��2�P��ԛ�b���s�Pp�h����퇺߹N�A�*���29�u7�q�$� ��R����R9GE�c��6Hv!�ب����j<�'���a�b�>�\��'�� ��IB`�U��:�KƳ��["��d饤 8�x_(i��4H���B�=�5' e�ۍ��J�~�-�ū�C�u�I�n`t&�����K�k�6䷏FFU�%���R|eհC��v��7���?�e�=�Ƭ�qjr	��l�ϰ��{�]
��E��[I��;+�,y�@����"�b���a���OP���m^�m��Z֛u9|��|�z�]+tt�����H���=k�����+���V72��dO�z{T{�T�;�3��
�/͊���Ď���LM���~����߼���I�<�f$o���L�h}��L�?0cSD�w�V��"�r��X;}7�T��hhF���[�G��Mo�#��ܮ��0��W�qf�<��� 0X����k"	_��K���b�c��x�H76�����՟��#�aQ[�9� ��C���A�:mo*�U'xf����ֻc�����\����R ����]�4��{�]��h��)s�$|usʅ_g��Q]YZ'�����I��m4N�2���4����N�$�s0����/7PX7��$����m��`8E���&��H��*Ȕh$�م��&�r�����@���������1_'Өl�6R.��0TDKZ�K�g�E�������S�������j�4���r���Ep���N��Z��"Ɉ���UiR��J-J�"���t�F�Vr��"�$��z�/:�V�JU����L�ȇ1�� ��
�w6�1C]����Z�^3}�m߰��R�j��U�W�<��I�?�_��Pa��^5���Ws��ӆi����Rx%�/���5%����Q�dl�u�o����nC`���z������S�g�HjV�1h�����Ί'ǳ�B:��T灉�J�}�9fA;�]·�d��y��䗰n�J_�2��3��<�85�LI2e�����	�7�E�P���v$_H@~��5H ��1��r~�b��j2ɿ�VzEJŶ:E���{�G��]ݼs�(NUO,)�;��4Ǽ�)x����5�����c����m���K�P22v���ZLת�r�!��6 ^m�Z��RR!FG6�#�J(��>
2���#����)w�c��˞�۹�@�4W�q�� ��wdG�p4��͛�'u��<T1-����6����2�L�@Q��I�hM+1wg�Y�
�G{K�3�MYqF�@��
=�����t����(���S�� k8F��]�Y>*�-���P[�K�V�@tʄo.J<"1�bytF�6��r�a�c�س�Pi̼���03�p�����?Y'��p=���|�O��?���^�c�;@3�?�?�.�)���?$�;/�b����h�5!`Ţ�_��IX�W160�$z&��7���a�l/��d.O�0�p��SB �j�d�䅭��yod�ld^ ��׉��t@��2np�&�|o\^�O(F~l�r��`S39�n�;>~-}�F|�c`�YoI2�w���1��B�kN�Lt5ļ�Z6hט�&R����?4c�s8��Q�8�x,lz���]��[��hD#	;Q�èj��jh�16��e��$=&pYfa�"��1i�:��i�js�_�a�l����U����ϡ������wqc�&�G��_"�eTt�����v���eL�����
��W�g�����R�p�+���>��J���0�n�n�����M�m�
6�nhc���WJmY�)����_9���N�j6q�kA0��>ͻ�}�#������lj"M�/�x<Ë��ɑ6��YlX|�t�Ɇ�腋��+h�YR����^����U�*MVS�P4�c���G�wH(�w�q�0L�)[H $��fVU�J��о&6�I^/F�|.�Oey5���������+e��8Ar=��<Dklqs�nk��%�5��;���� a�L�L*iB{��;S�;w��.N1�́!q�q��{�Y����T4����W7����	e^���yY�WoA��:��F�yR.�&-���@E�k+��	���G@5+��l@#"Sq�8+%D�t|됭�h�&�,�¼3���G�p	�����4N=�.�6)�g�_�-{�d�;^@����{8S�=T[��<Z�8��8@k~�̋���V����B�Lz��%~Y���%Y�W��"�	rs����nŻ��� �����,ʃ�5ŕH
/"=�wx��QLe(eJ~��+}�֌��ai�JI���]X�k��J An�8��q!Tu��U�(Y3�惡�;�g�piw��+)^W#��8:'�'v��:�n��Y���u�}j���^~H�D헅�ᐕZ�&�]�J�Ƭ�Z���/�Ԭ9�(��"�H�sU��CX=0i<�^m�ܶ���S�lP�D%"/k��jk�9`�9m�� �d7�g/�~��.$d��i���}��*�Y܆�Ȗ�;"yKÒ#�Ť@�hcn��X�c4�@�e
Enf^.5�X��w��k��G�3���uq|���X$�_�b.%��l3X*^�qPP�Me��y��|	 0������\]��o0�]݊~ ������b�"�I��'G6_@w!�8�7(�n��5dC��m��Q��"Hx*�V������������(սX�k/�',�I�`�>�b~�X�V���������$�I#
���Xk�ORޯ�gc��G�~���5-M�z���J�H����փ��y����;�-W�Yc�P��v�'R�b�� ,B �⃩}\r���������d�!߈��]� �d��on�W���Y+��1�et�:18�/i�g��H:�*D[S�e�B����U�}x�P�| �wڜ�{��R�="�&��0>��iL���}��$cԥ�wF�kwoy��/������^�|?��j��3aM����'(��1P��(�!,r�OU^{h�"�[�X�3/�����{���ExgK�Thڦ�xvU��!�K��HV"���ewLo� ��/'��$E��Ą�F7����Uؾ��k�9��$�5���h�ޚ��E��A���'���8!�%Fq�AE�D���ƌ�Q���Ԙ> '���۽��l]zQ�[�E�Q�By��eB�C�"�R��rIb��2��#
*r��7�M����]��!hh��fgn�iʈ�n^z�#�z�g�#,O�c�s��&(u9�]�����|��T�W���wj�|M�m{k=E8K ��2�B�^pAF���ǎWzU��ONt���i�c�'_�*�Y��i}7R���*���k=;{.`\�7ғ�
��㮹��K��d�QM�OJ�������u����O�7��w�?�1�Xvt�1 /pkMQ�Os;ЎL`���d�Q�Fkǐ�l��4�����0Wl��&$�
D5�߆��Ⱥ�.�խcW'�s�j���x�w���0Cbt{t9̳ɲs���zl��X�Hv�ɀ�@:ys5��2�F#~]2X�JΚ��S�d/i�.xgdz[!z�2�E�h7y�˯�ɭ��l�y\R��ȓ����A���J��?_�����c�EL�8'*M�w�'xK�TK�߯�w:�D`���6�!l�	X��4cK�'aaV+@@���N��*uV�}�m�7�p=�#6=��`o�6E���u'U�V��#_s"q�Pd�j��&��6iB�����TśY��)�W�d�(���R	��R�l��/��t�S�釧��oB����O��+Ⱥ�����~g��]c�t��MS��?��T����_����5k�yX�K�I����+�~@��ӵ�����5^��j��z)!����"�@�煂������ʱ��#��'ʀG�u�<{Q��I	���g�~Bg1�V����g�0��y���X;�����F��l��nh��
-�c�r���d�b�9b$?���@s���.$s(=��jÝ�+7{n���#�3�硁ɯ��I|Nog�tJavRE3��7�aD�P16y}m��D��[�	Ѫ︄�i��2f�k�J���a��S]��ΪD��y��㹞j�6I�b���}k�����ϊ���K������'�G�7�ZܔpI�r�\ɇq�;�Bq���T�ʜ�*h�|A�� FQ��Y��+�;�p�mc����/�D����)��#�L�p�]x����7k��=�v��b1x�[~�k��ik��&���������}]�Z(d�ڶY�W������)w|�X���
��_z���J��.n�����B%�B�qq�R��E���4�p#g`�t%I��{�m�q�U����]L�Ii4$ӌ�,��0�j$�-3����
^<eP 6��}���opESJ���i��V��as�i &K�n ��ނs�N�łW�]h��� ��,W��5l�����o�>1�1aKI�@����w�ء:�7/7��~��hN2(4n7�F�^�Ö?�d�+�0���8F��&�Jg�Yĝ-q �|�2�ێ�OXX�JT�_�쟖�Jb�E�����{��p�N\��\�����j�C��G0��������.�nf��)L�M$��4��u�2^�C Ie8[m ��}ȧV8���s�B����y�-槔]��̝�+�Z�`�T������kS��ӟ�mһ���H����i�P'�˧˱��[u���Zg4d�$�*����B�ӱ�vX=��"uV���V��ob����%�Q�lwV�
�,>f��#�]��Га�D��C[��)���;}_��/��R�دri�4|�Ysm\�K����ȋ�M���b�� �T���s����f5�M��)|G{���Ư��V���Ӟ)ȑ.�Cmp�V1����\��s�3��wy�^@'x�!hڤv�'�j��6hۚC[Qvz#N0��Z6 �e�	]��2�޼J�������1�$bQ�m���f5���-$M���e��Lp��yBy��H�akǑ�25M:������A�|X�+��4��G��i�wpi�1F�.rv9�����N�3��6����wd��;�;e�K��n�/�,V˦~��"{����*;ͦ��c��!I`�*`[u������^���/��y�0R�3hz� �����J���;J��I��e�bZM��$;�C��ū��zC�5��CHJ�4�Ї�&ۏd�II���<�7N��0�y�чi��e�Tܶ2+$�>d&B�V�d �Y��i�-�Ӏ/��F{��/C���M����^hx��VU`&[i?v���?s��#��¡�ƚ���Z[*�Y��3#��޹�:_7f��j�Ah�m�o�w3X�LT��k��E=���� RC�M�\��	�bN�Jt��X�������=�ˉ�f%�P΂x_S�t�v�}Փ���f�ԙ�ՁF`q�t�����xe2cm�d�b�m$u$��o�Y��aR�A{x�G�9�tW��޾�B��)!]z��[����®�ltP��m>~չ0|�~��O�a�v[DG��H�J9�X��ӥ���Nn�e�n��S����\������Q�U'^y���_��64�2h�Ɔ�0�+g��P�=�J7�����T
��m;�HVfA��s��K�hmz~}�D|s9	����b<��!�w�y`���*9(���ffD��Ґ�0?%)��J�h�ֵ�y���K��?C�\Gσs����d]@a�K��}Q��B��$vS'��RW�`J����'bku��[�tv7�^���iy��c�����47,{�>���~/�}2�B����LT�����`H�G�?]䭾/1��h�)λT�¦}r�\0	�C���|@���{[�f�0G�QG�+ ��懝��&�APL�(ᶤ�"��Ì�/��5�4I�@cHC�6��y^�"Z�A/���i�� {<�P �q�~9y��C���Dp ��RM�Iy�[;z �j�����WJ�ak��Om �}��ۏ-��V(�v��I`;K/� ����B��E��_��y�'��)�`z��>�^�
f������������<��g� ��v��X��D�/x�v���0~�A���V�nM.����[2���lǰ;mE�G&�֐�B"��V^B��O�+���%���Rpǎ��Rw��LB"���$�� {l���9�� =.��{3�f�f\k¬����c����c3��Ɠx���O_^�1��2����1(B��C�Gk�P�Ɩ����6�T�W��Ϡ��G�$��Lyf�4̛�`� �９W�xs�81�%�&a�{�^��͘�#)���2��V�bҘ c�$�9;}(��i\2��Ѕ�$����I�O[�;cX�����k»��D��$3	A�
��i$5`�����pzL�P6�FkdA=���� G1�y������=�Q�r�M��?"Z���%@�GϤ;ZւXF��"�z�>&S��r]�;ύhU�Fi��{�I��|Y<��|�X�6�y9�����6�f�ȂyQ�{�ė���YDrފ��@��Ӯ�Np�.s���4��u�fb�VFki��"ff���8��t�踚#W�.�L���M:�%���zn����z�qMڕ1����3{
�7�!iͻ���g4� GD�)nW|�������xᛵ��`��Lq���F"����M;�"y���ʧh��^L�3Q�&��u��Z0	�M�tp�	�NfQX-�P������O �@�&}�~��-h折� �a{A���,�2__��h�4<��l�b�r�M���x\�!��+��K~���t���Q�O��7J���b18&�a��CԨ���	m��)�Jա����Y��uE�]9>}�c~H�S5N�����s��-�@����*�G�p�me�f�z�&�"�S�)��p�zx��]ʭ���\�DR���T��}���f\�����^���t.:~U/&J�z7g���OJ��y��?��E���:��^@*ѝ<H��5�j	�C&�Uũ���\���Ӂ������\P�܈i���%���!�	��%��k��	�N�����'j��!Z�~�Q�z�b�r2�և��'{xV��K�}D'T��<H?�"_���b��g�K��{k-
�˝�{�\���h+@����A���'�@�Z�~2�8�Ӊ����0:�'~���w�z�L�Z6:��A?~��e�~�:����6Fn;iY�\nkN	���ۤ�s�|��DV�����`����3|ҟ�H�GZ��TqM
 ��C�*�elk��&������d����N���~��${��Op��ϐ�Y+so�^笊:g��a�f���n˖��W�����W�z��u���኎�CS�	��J U�ˑك]dו-%a��J��ϞA�D��]N��poG�Q"�*��$V��6��4i�l������j$�����������_.*�#V��~�
^`��'���A����&e�/��ʢqD�{��JО+�
��Y����?�ͣ�r��������#`:ܱg�z-k�_丹��5++�q�%}i�o��xt!�;�M�c�����~�P��-�P]>��چG���i�&�8��%�����y����/4o8�
똫���7��"��xx�C�'mr	'�]t��ڻ�u.��Z�:�C�Ҡ��X�kB�L����M��Oo\ivN��Ϟ�@������8��8��_�_h�i��"J�i"�F�n�6j�Y�D�M8#m8䣓 �����9���$U��\+b�5̈Z�-�A��t��킒]�]O���H(�d\�����>�����5�"	������q�������@`�A��������V$2�x�_�d^|��#��i�tfoչ���Ss�-mũ�U��y�c�d�	���E�l~�`�5�}▧�vW�}F���7�X	��o�I�j��T����_��T�ѵ�e��/`��YgA��O�"B�~��Uyƻ�Ś��ȴr���?����ĀƟ��܄<�#&S�4*a�AS�toP���7U|���tLH3�2��9���v���br4�*a�d'�'�R��ٚ
��fGc]:�%'ucS��7@�-ddv�?�}@z2���5�hnE}�����a����F����g���k�����>ȮA����$�3�]�8>^gΟ*��KElW1#ˀ�߹�J���.wq���l�bȿT9�|:!2�S���e0;��7��A�8=&���>�I�ړ�Jd�!R�s��@2��ZL��:������O�<_����qڨb��+&��KD�ڑ�;
�h�+!��5-����c,��zU�%��MU>��|C��Z����AɺB	:��ցw�!9"�OD)�$���H+�3q�\Tq�DĀz�ap��n�DGfO<-�`X9�=��?��[_��;z��G�hCL�eQF4��Q-�K�j�ϋ��\�&���ܛ�t�:����TL�<?Y�g�qF�,@e,(-��3�������v����-��u��]_L.�E��\�*��W2�X��O���,YRN�y�흭U|�kc����'?�@��_+|ĮY�40��ir ȁ��$��(q�OŶs���=b%݄�b����O����Q⸳���V�T����ĸU���	���W�O����n�8�`L�F={v��_�L���.:.��L�T��{���PaX�J�%��O,�Åڙ�z��ù� @{q��:r*4DH^����]�>=�F�7�[
�������g ă�{9Q4���v�tILф0�sX7�[R'��SAS�����S�<��zD���y�z ��;�CP�xb:':��%ˤ�d�L�����`6:���7���jj���cל��Bzs�!��8�RL
&���3�TP����΃]tPk�Z{�,���z��?=�J�{;�%pA�w����Q���������j�'�㮰ϤzY�%e:|���.9MWc*�o�Z���X�[6\{9��5��Į�-�I[k��Ť�'1��Ӂ���u)���$Q�9��YAmb��G�>¿ j�i�&0R�FP���-.,�����@	G!���.�uZ�~��k��Ny�Tc��O�dk�W��c:����2�\�d�i�e7�����M�Y��8�BY]�y�W�3pb��B]�}��]7<ն�?p��/sg��r�RiZ5/�6����m0 8����p����"�H:�LP��L��E8�`%FQ���<����ʘ�	�����w11���8��^��j5a!��
�=:G&�o����N��n�Ra��1��9�����bq�-%��}��N�s���<p~N��{���ՈM	������z�{�h\8،�"�L�+'o�#��py�_p�fGo�~�T�j�����O�M:Mg��x� m0)�u����Qh]rL�՝�K2!S.��o>G�S�l���b�.`
���a�<�L�[(RI�(f]�"�d�}�*��"�(}�خ�e��踖Z�{�k�z�B��^��x�n���"8��?T���\P6%L�̓�UZ����k��KkGg�s��I�[��������o�u2��T�g�~��	@�F�����dg�<�)�z��{�d�$6��@\��1�%�n�A[��FN��^�N�	q�Ga�򞶵�V�ƑN@��e��Qx,y�HY�1Y�xN7}�=$mk���u��x۫-�$�5�}A���
�coF�����.Df_���Y!Pr��<����b��zd+e~u�:��JD�|�T �~�� Lc�#Mud^�� ��v*La=.�fqXM��~Ͼ��E�`��/+�K>���\-'���k�ŋ�[_�.��\v��"w��hE�#�O,Ө��oC*IAЉ*Gf6�J3����ާ�I��B�T/ b�eÄ�vs�K��蹅��y�>��îޤ���x
�ĝ�@��u���mCu_�y݈�lߢ�)��ãF�Z��{�hN��3�/�+�.�Kpv��H/�3�h3��M!�;���L�����]�jFե�b��� d�:K�Ӣ�F��;u�B�p+3?��}��6��Q
U�D��~���)��L�|\>���I4���ORc@f�+��|�ϑ�į�	�4o�bϤ��V���;��u��|:+Y�y3�?�9������H;����������Iݴ���ΐF��;��K�P�x�O�r��1=PW ���,_" �0S��8�^r[���g6�뮠��	����|9��Ţ��A�r3̰��9��L/ f�[	�Ԧ��ENJ��������ɠ�Լ0ѯME�%��<�G�"(�ko�������j�(�"m�[/=?�{iT�K� �gN	�3կd�A���To,�*�����YAh��j/� �	I<�Z4� תh�X���'hr�1|�sY,��B �-ɔ�Ƽ�5\��^BW=HZ���D�&�Ͻ6�D�Ĉ�p��Rn'�y/���������A�7)�1l��x"`a�$QQ�����ij0@�� �ڗ;��L-3����7[e' �R`���̥��ܥj����ƅ�L<��W0���gd��e�o�OI�<u�#�C"xWݴ��?M�w����M9���?=Q�[�V�MK��9�3�9Ƴ ���æ�g����[	'8f���呀�[Kg%�n� u��/���l4/�O�*����m��Ù�`I����q�%���	k&;ᐠ����6�³B�;����w�W�a[����u�{��Y\�o]2��d��-�[B@���8��+�9Rqg2Kqf��;�u��s�'x}5�R�RD�O�80���	
h;8��kF�ŏ�����N
��G�/���]�۰s�9����L*����_��������2��-'3�jS9�}{qf2�7|KE�f���:Yo��N�CaZ�������dՈ�VC������ɦ�ɜ�f?i������x=˱�`\���*�ܚv?�\�R����ԑ���F �k7r]�vv6=� {�{�p#�_�D�xs.9��b��^r�$�?-��k*ԝr�ڀ�P���y9׈��4�������)\7�l�Ew�ĆtEe#T�c8ǰ`9%1=���� ͸/ \Yp �^�¦�@�`~ީ�a��-/DF����흂���ǒ���C�U��4SN���1����g��K�-�Կ�e T�=���Z �7V���G�Df��l9�R	���J7	�}1��Q��S.��Y�x��>����c��˸�_㩽��6���sM�j��Q^R�2Y2�a������(����Zs%��ї�U�s�#�4�3�1׼%m)����~s�=��K�S��@yR�J��!�Z�Y@�1;R�&�w��w��m�7BN��55���@��������՝���"@���q�^ؘ
`�C ������I�!=�s%/���*Z/O#�_��ԕ�J	�oW��%�@�-�Q�vvF�މ�����/��c$}���=v�#�[S2�q���i���&0�[BcB�PZ��n)�����f�ϫ�O-������>v�ا�k`�`|���I/��?�+U ?�!� �D�)??e�Ԁ����#j�p>6�Xk1Q6��{�dr���i2��ߍe�����u�,^x�z13��5����@Տ�Tr"�;��/�+h�D.�l��Kw�����n��,V��`$
�.��6��)n�G�(m����SK�8`A�縹1aB��\p�Ui��(��U��X��)TD:����!���}9!��_US�,|h�[CP1���c�̚I�Ӑ��M3-N��D$�.	'�
rE��"��v ز� �rZƼٛ���mbk�o����\�C�9S*BifL1�#�,���E��k01�/��@F	<����ܛZ�8�s)C�6~�t��L1�M��a�M�ł;B�d{}[���~���\K �S��y�����b��
�n��P.���+�t��b2"�io����_Ms'Eҥ ʹ��c��d��U3wڼi�_�g´d�4�ĀPr������".*7��{�.33�<S�c?;�v8��:E9_`9/��T;�+{�<��@�g"�#,c����[�=P���~��f���&C�n*]��o��@p��e�I�����-5��{Q�6Ԧ��%�9���_�i�$3`Di�};ԢUz��yeO��f����,���!�\�8$��$ �̩0Tƨ~�u6B��A���#����ŰT��OW�
q�n܋\g��I-�~>������i(���^��l��l�..��Y��N�8�`��I�X�/����& ;o,W��	�:+��3,(r�v���}���f�]���?2N���͵`m�ƛ�^�R���)%�>k0^l�� 꼫.�}�������t����Ԍ�dXho��ƍB��!�d��8s�yRC���Qy�HQ�*���V�~M6�"Qv���I��Z�'����Y�j�f�ē8�N������pw'�v�y�k�]�ب�@�Q�&�S�1Ǭ�&7ht���N��r��V���Nr�#�Y�u���H�~�G���Ry���Ȁ��3�8\��6��hO�8��U�$�.���X{6#p$R��e��ܵZ{�t�&b��d[��%����ż 7vQ�:�ξu���fc�Ϩf�y���j�W�z�7�Ǽ>�ݤ��b��N���0�!��c��c���M�_�A/��V��g�����`Dw�I���%K|"��j��tKN"�s�D���ՂO��	p�h9�����ev2'��P%D���	�`>	,X�}���]�^*�]�q���E$�����zU@�ۡ^�(�̹^����il������
�c71��s���,/�6&���:Ƕ�ΚH�;��읯�a����|�T<���w��B2�da�?���ϫ�����A@���ϟ|��2�Г���VN:n�r�q��e1y:�Xˢ�
p���R ��
 K�ici)XeK���E�bR�r�brB�h�O��9�Ԁb���%�,d�ᾖ�;�W?2/�����e,jn����]X!�BB.���NցY�����Iw�{tRغ�+кr�
���+���yQyc[8`�;�|�!Sߡ� i&�� R��C�QË�u����{�ٴq�|�t,�T�,�Մ�����`��f
��P\T����L�s����MDZ�`ڿr*�H��.b=�(�YV�z�la�i �J�7/#
��B]槩}���M�K�~�қ���T�C�Y�|��}N�䝧���S�Z.=�8O�F��9��5T�&�)��{M ���^�3�Kw��!�+�±SU�S�#�4rot>[��
���Kr��z)���#�9���iM�U���?�䮢��D���5�p��]�Mp�Qgb�;}.iuEŠ?�s�5��%G_4�;�?�&[��HZ���G
�i�=g�R%d��fߋ���D����e�茉2�nR�)j1_V�jm����<� �������|Ȍ���~�2����ȅ��q����O��*h>���F��Mp1�/l(��ɿO@�w�8�?ᴕ���D:r��N�Hܹ����z+]������Xϡ�9��>��}���z�l�h?�Gvdp���v�?L-�2�Ws�},>RZ�z��W^��J�J���i�T��"�2�R��y����	��T9�ڄ.�~m,�m��{����	Mi�h1�K�*�L謥D�լV%=`�U��"7ZD6��=��Ϣ=V��A��a��\K������pW�4��U"��T��f�C����`f6�W���J�PM���g?d�p����{Zț~v0@�~���e����� �W�Q�+r����z>jh�V3�'#���&_�D���'l\$<a��1^��%��j-��b�:�lVB�q�M�q�MZ��i��(�*[��|�����,3��ح>�*��,�$6����>�~E,k���,nrKC,gF�8~r��9�vBg��s5�^��y��^_��^2�q���"�8�<��=qH�5���*&���]���&�F�^ڕIt���c�Pȑߒ2�`
);�ڦ�l��%����L���@�ƻ��k���{��)�^웓�\�����=��"�r�wu9#��KQ!��O���ݣz�ݦ��0g��:��E�} s���>�5�q$[1�;d 5�#�S�*�X��̿�-���|@����%��T�l�'�.׎�7�!O�]�sU�V�5۾?c�7�f\�`F�Qy�E�'�϶�=����8)Y̅��K;�?z*��qr�xOF-��9oȸ��ť��[%XqR �^�G�2�u��Q�Y� �\��I^Y�0��>H�������S�`&u��.����몄��sЋ��	ѡ�U�?�w�C��;����i��x@N���a6nƐ��=ax�]~���Ie�FivӸ׺�<��xj�{b�!˙��r/�;}�IJ�~�5PF�n;�(�b7��ey�H�1�w��t�TEؓ�������P��:wϗ��˜F�Uxp�5�J_��t�Ǐ$3ދdB�5��`ߛ�CN8��O��F�i��Fr'��2NT�M�����8�S�SٖN��12 (Z�����4T���^Ɯ����K�oY��F���n|X��+�QZ)��lX#��(����m�^��	��).<}�� 7��I�G��lc���ϲ@'ʱ|Pa�b���pd�{����  LE��E�����"Yy��H��GZ�t"`��4σ��Hos���R�?g�2�F.	؝���L^q.Ѣ������R%ѿe��)W��� U�r��G�,T��$�B���)�h�u�Q§̅������!�8��"�\������K��~y�;�1��a�����AJ�C���V��pO3d�I��R��8w�U���]�+YE��ڨVJ�߱�KXUfL�0�T��6k93v�|Z�0�'�|j�+V��5�ԟ{���Ddy ���5��'Y��'%��Mϣ������,�en@r����&{_i�A2𧐖����)2�"�4cDTqM��Я N%�r<zWP*)v)%On9iv���B�,�윻��6-'��G��N��"�	���ɒY<SRC<�f5����
�f���b��2L,���,N�Gd��LY`PL����+�͕R���B2/WK��A;�ͪW}�(X&���~i�N̓������Tu填<��g�h��o��BK����o��Z�]/�߈���G�=�\z��� �j�6��?��}�������"ld��T��C>�>�s�����4���^L��O��5z-��BϵD!Ϛ!�^��_!vR��O�����$��2���V���{T(��U�V�cw�c�%�Y����T����2\B��$��aDJ����$��4��+<tbv���Q�����`K��T<�L� ���zf���V}�C�s�?g^�R�3o����ɀA���tk��`)����O��'���]��j����)���j����R�Gctإ���ܦ�QSWP�eJZ���?ög�&-�v��ΥN˿�ǴHօ����D�ă��2�$s�hk!�6ыc%3t�R�-,UR{<��n�w�.��j�����d+��	Al�8�ӓy*=Y��^dw��P��y�} T�t���������?��&�2U~����o/k6n�y9��c�Q�,LM��R�"%�T��@���t7����1�p!�1Mu�jJ�Efa��;��r7���jx�&�LYD<�bn��P�]@��>� I-��.sPi���^��VޠJ(���'��q0?�k�-t�٥~3�Nt��� #n�N���\F�3 a�7dD%�Q�W�ӽ��6�B6�����i��(̟�rO!��� �������8�R�V���;^:�3bW>�|��[ן}P��-���x��HMy��i��څ���2�jk'�?�r�$�2J:Y��^�_\�^��c'ϵ��(pa��������~Zŗc�4�Dr#�� ;W�H�����X�����F�/�m�'�`#���L�����h��+o����g��ڟG�����i^��M���\�n��wL���q��4����6�iP͠z|���&��Bp�;�$*�x�쎣%������Pu��j��t�0�N�?�����;(u���'X�AT~�o�i�Ʉ^�g������aĐ�5�iq����NP��x�P�L߅��~P�Å�V� �!�hR�!��6W�-Ϛ�+�H��N_	L8-�L��� �zE���� �/`ۦfQ�z��!��e}?!�p8�3�U�N%��'�P�����ɋ�C��!�x���M+k�`�/� @��8�{McżlN(5�͵"��;([��@4d���|O�!B�0����*�;��m�9f����T>�����W��MoU�d*�?2��2b�ʅ���vb5XE��m�OI�b�M��y�gZ���S�6��)��:i{'�ݘq�h����x�%{q}�����U���?rr�,rd��H%Q�p���G�_֎�]����lзL��^ʢ��Ih�aN�.������ )eE&���+zꑳ������ej�I�|]>�{4�� ~E-�|H1�8�'�S~`8�M:BP��Pd�����$�8�c�=��[BO�,�㤴g(9Y��!p*TW�(��+Y�{i�p��l�V>�h�-\pc!�N.�3�\��5J8�ָF��p]�S4yy�
f���
FfYŨ�����G
8#�wǄ΢�*{b��B�E�����Y؀��6;�ڤ�F|!˪����N��� PL�*Rdr��H�:_���Xa�pc�H>-)�g2̋:�jZ1�����zRn֌\�zť2��o9�h��Xt=��>��0�,?h�dA!9�.�M~���
�=Uzl��c����q9��J��nk�V�w��B�2.���H�C���_�
�=�5�Ǘ/�"n�4l�w}�2�����qi&����ɕopƠ��6����4��YҸ5:��N/(U����?��T�h_����� �)>�X��	ϭI�T���wD�	�tUb�0e���mL ~�(�P[���^P�g����9ͅ�����-�aZ�����ѽ0�7[��𿡩-��t��t���gc�k-�#7#/�3m:�j��I_���]��	)7��Z"74/+���x�<FӋ1��a�ف�3{�B1�p�p�)lWO-9�B�^�uZl��������Vq>��.Т���)S7�z�x�hXO_ϱ4�@����w�&��k�s%�����?s�]5�}�s�x0��)�o"3x� �h��D�|�?�y��}!�m�"�ݱ�Ä�spWR�Ռ����ŵ����+�:�� �y����  �rF��Ay���  |�,.��M���af�R�ZAl]��ҩm�H�
�A����lA��$��d%A��B�䒛������0�L(�'t�ly��/Ɂ���ӟ�P}��`���h�&�ᓌYʆ��mTǻ�9%���(Ø��	�4i��5��
]Y+�F�wY�͌�D�S��O���C	���섨B��������J��u�y��8�<���չX� �[����d��%�k��3�F2=��)��MKb��bB�Ӿ�
��d��2tR��hs�޹�<�ۨl�?�⸖E$5�1��[��v�߇V~��Wd�:0d���O��֍RR�sjNe��.�;�u�zsE��q#	׃�PD��]g�O4��Z�IH����^�=#3�7g�/����y���M�E���AȲ.	����38�C�m�h�
wHѻE����M���Ł�@,t�MU"L{~���˼��c�8����*v(��i�D���P�����c7�d�e���ӥH��m�>[���
�s�Z���٢��&��|pe	��T8��m�#W=����_���34\7��f8*J�iޣlc��?�/�3��Z�6�k�d���OJ3��������2]*Q���c��;ZP^w�ʹ7�Q��)�f�
� w2��B��P�g��lcc�L	����s4[=N��b\���'��e��ix��A�C���ᯢ�!��d ~�:{���b#s�a^ŹT�P�����<���'�A~Re�2�YU��Y!UA��1�e�(����+�ӆ5��$����]���_��1"�<�Tn����-
{��S!���+��t:q�u@�pt~n J��:��JMR�j�� �SҜ�p�p_/헆(�}�}͢�'���Y(Bmb���-w�a�����F�,f[4�hƢ!.d�l���Y:�zS��6����
<��O�k��A&q�j�>j5ʐ�^�w[hr
��
\��S��s/�^3R���b5�d�{��FKmZ�0;�ʹ�lE$�5͗q��\gr/�� f�+��͚5r�6�9`��J'V��`h���&����Iv8�O�a�ѽ? Jdr ����"ޚ��_Hԧ�2b�,VL]��K������R���z(iz�<�R�Q�Ang�xO_��%^�-O�/�[��|�I(a�6M ���AС�'B��ܘ�������:�JR5�����
�Vڈ��`�o�j,{O�� ��C m�5�hȦ���H?�{'�Ko�SIk���f(� ��ŭڦl8��@:��Ol���h��[����z)�v��Y�S�أ�}MR��@a	rO���b��,����.]���ڵ.裡Ѕ��z�Eq���t��*-��Rg9�����f���U�7-̙X�q�ׅ
0�-s^��_�_"��:]<?��8KQ��r�$ҡ?�|9IB-�a7���F�;�7�c�<L�`�L����}SGi�t%��$�;jzz7���I#�`R�_�NYA�S�sÁ��%�2B�@^�h��|���I�����ux-$iϖqV��&���/�VE��;Ə"j~�7���WA�7�F[�Nf�*��2p��ǚē8Ț��vZ��hZiA�xP�k�=�n�9��K1��F݆?��\��˘��9����%�
�'YM�+�[IG +�t�O��Rz��:۞\o��qi���f<A@�-���"�A�*W�`Ǐ{�M��`{���Sj��!��=@� Te��9dڼe�[�Z<��hpC�;g��1��FF�Z�" `�
�ug:Gy���8CJKT���准��BU`@��s��e.�S�.��`���PGT��
�`�(B�v�xaQ���<:�m[�P��p�5}�C�Q���ɘ����J@�_Y�������cS�}����秋zm3+��ǉ�:������٘�d�Gs0hg��*�t8JD��Yt�v ��l��(����Z�A+%�r��$D(5�k�<�+��%CXc�v@٨�b��7�&PP�i5X�� ����]؁�L�S�%[�/ٻ^&�3(����4�rZ�Q}��;>���L��[,\ n�c����5�S=�����R�5g�E.��ҭ��rE!�Q�8��U�:���B�0ve�b���(�E�Q�c�0R|֫-H���i��:�W/6ҷ��@;�Gc3tK��HcC�!cM��m�aG�AX�5'��(0L,k���Y�tຈ9{�.�oU��m��}.�!K�@6b�#�Hr8',�Ŗ��G;z�+B@Q9�=}��7<Y��v�B�% ��k��8�?Ι��Z�﹢s�Pg�B�R<�2ubohS�.��ۢ�4�������oZ5�9��������NE�W�>����."?��~V����^?���-�6e�u�����[��t�5a��H��ͱJ@���\D��V#8?	,h���9�
����k��!�]��B�ۖہ���d���H3ֳo1M��)�ȇw ��&�;��wښ���d�ޮt�`�T?���&�}�	wWO>��n;�0�\jD`_�"�z\��n�8�WSVRf��<!lo�Xt�_괯��l0�̃:�+ޭ�&Gj�����g�j�8��}!(^�bkgCa��_��2�Kc��	���]�(������ �iܚD0�{�EG��8�qH��c�2HMd�h��،n�d,�6��!��%���:�����3��ʐ�uU��Qt�Rz[��z��q�G�gL�<���|�&����QG��1g $����L��_�tҐ���8qc$.����q�P��|DzE��l�ز,�ܐ(�l�l�a��K�L>�S�Z����'aD��l������,����5O�z�"��(j O�@)��)��)H���j�f�?P���aj���Z�I��]ACI-RJ�f-�\; �qW,�'�-ci��<7�P_}�Z~y��\���H�y�u��?�6$�~Ƚ�~�^q�ܬ�V4�\W[sĖ'uH,�>��8]-�W����w�e1ٺ�L;�u�=t��U��u����>]�l���p (� ��[��X�D^Nel��G3߱�W�zF�a��lżA�^aoP��))��2
O�V��B>'C����*ԙ2u�)\��z"���c������"��`�]�\Z���>��h��2!t?��L:&���u}|�Q>��e�L�4BS���}gL_�Pj51�CQw]Pw��";0}�s��6�1��)�������k<�K��Z<:������ѯ��<l��F��$�MupW}�f��7�8x7��g�����>�eqz�B�T��@��$����{�'��p0�{b��˪�$�����Fz5��k��{��~��Q��[�%
�p���6��Fc�k(��5���Ӭ4��|����;��6��\������3�x��9c�4��8��.-�R�Q��)?
����]W���,��@eQ��4�����Wni{f|R]9�@ 19]��}U�a�V�t��� 22w���(+���jv�Ų&�jz�sTkh;tS�^���י���_R��m�8�=L�r��\4�nq?$jq����LPѻ�1(�)�Er�Z����^����J���.�_:��	�%#{K��S 7���t�� 2s��C��:��EkbQ�M��o�WA�r��m9�%s}�A+[R�g~"�:ۥ��\,������L3���R�8��� v΁�������q��������e������֨d9F���3��[�QmLϘ�#ޑՇT#
��n)�۠�!����7��c���Ϣ?Q�כ�ݖmj}��D_j�����}!M� Fx��`����C=&�Q����|���,5r�Ohr��y�+o��hB���{W�m�I��Z\W��bk�[u���]�1���V�v(���R�6�u%�����X��`�6���[��;� ��!�0�O��~|��w�n���kw���v�A�Z�{"3��6������q���t����m��%�C?��?��4��\L��Bü��	�cP��t�GM^z�F�o��|G�F�1�63(�	�4�iU����s�ӧ�g����X9n��\�B������e����3������qKRp_D@���t�Ԙd�(H�<�h���Z�*,�&�,V�W9X؄�p�ʉ�4>-������o#��AG	�.27)I]\�� �sDʤ@�aoh�KP	���X�N�Vc�G������}0{�������,W���i	�����xM����8�#�b�Y9�Si�ҡi�}n>C�H�b�퇆�Fh�W۹�^�Hx�� �b�#G���^f�@r���μ,J�7�D?+�/!�����.�����]�a�z��}F6� �hK(�N�Z G�%�zZU�j�H��f����(�l;�HS��Z�F���3t\d�ѓ�?�{�$�d��:}�\HMF+��PA6���0\�{�V�N���]�{�e˯&�r�'a��ٝ��Ild��K��w��֮l��V�6ىj~B6 ��;Av�}d��I�NqӹU
�����*�š���ג����z
�(VBU�l��v�����|J@�!f�KJ�-U�U��D04��G�JXIt��s���/�A	�*�=5�vWF�����<���#�R'����C� �"x�r��0G.�P�t�x�t�����V^�D�� &�n_P� #���~�9��MF�h�l��oEj�mTֽrI�@}E:�`t��ܷ=f�`����[��Ӱ��-�5�l��8Up^��>���-���e?Ш�Ɔ��I�|7:�u��l,Ft���W�"�M]*_<ʇ�r��R��^��61g��#���H�B|���%W�6M�}�W!07z�~���_/��������XA�;���/QJ�}ml`�e'6�Q�J��D�!�o�'z�=���[ԑo�\,j�TWW�9�����O�U$�N���}�{\H&�w=I#-��-[Q�W,e�6�~A�X3��� 	v_��a#��T�@HF�%��+��Ư�~֢؎mϨz��YY���BY`(/]zV�����˃�M�;��]�C0�c��ǥ��"/���UO�=q�>�L�=�.12\�I�b~�{^_�H�ބ�p�$pX��r9���lo�����nlڊ����$�թ��œ8�4V�UQk����~af�, Cn�������AuUŁ��
�cP�HH��s�jWtJX�|��ދ����*� %���=ZΦK��[�����FG�WWoǣ@�,RɎ
������bv�U��Dh8t���#`�;�"ı�e�L���$e'A�d��`�Y�Q���N��߱���U-���>
D3f`�_w�6��f�� W�C֪�r^�u���`�
�2G_���:a�_�FJM�X�zP"�{�X ���9%�B�ǲ϶
�ӫ���a���:q�*��s�3�s��)��0�	yr^��a�e����P~/r�E
ƽ����~7~_����Hj�-��;�.A2�[�~�������2?֙W�y���� h�a��7yt��0��Ë-���Ǿ�j����P<��\���u��9.`�����!�?�_J)��[��6�S�nm�2�W��fu��D C�0���85NS�@�@����\^��ʣ�v���4{gyk��ѹ�~T7[/�!��s��Qֻ;�$�kБo��\�O̷Ep��1e+����p�篅��^�V������4��z^_$����{mM�m�!�r�-{Q�n��MK�8s>�0��%ｚ��'��3�����x_\��ɉ���i�ݛ7C�$U!�t���r��Dr
s�A~�LnJ�?o��� ���^�<H�ޏ�?Vg:w�J�H��{"B͸d�1-�fq�r~�	�� �j��B�Z��x��H-$�=i �T|\4K��r�b8a	%�xL:���;�B������d�`���)�H�I OـY�"��(��冼��+����Q�>z�֛�>����q)����b�ޡ��4��[���iL�v���s��g2����BA�N�=>��r��t²(u�T����W������9
�� �d�ąT��RQT��i�T�!}]N�A�j��1���	��%_85q���Q�h�j�%A< �OKMg��l���p���T�y$�t��d�0ޫ����ЫކD�zj�W��>��1�½���w�BBHZ^Z�����A��2�z�����X�{i����R:�%;������U�c^���?f����x&
A�a�i	�"�T�/�:��n�#a:���#Ա/~�Bw#l��ψI�-Xƒ$�--�WgO�9��]2�|��g��	x��5�O{tM�f��L�!�	���g:�$�GP;�r��ǉn?�qR+��y���O�a��� ����Q=��!�C�c����)�N--Az��WA�1~�J2��[ln30��f�F̥A	���#n���܈IF��֦��fh��]'�k��:���L�A�,���i4w����`�.���7��'{��X�ue����LAU7.�D�V�L�n+����� �C�Q�c�b��c|u�r#$�}��i�T=��5#B����������������?�`fc�K`��.��t�n��#���\���Ҵ���@�>��:��v&�:�u�;�0L��L�ݮ��βX�(�`��?�G;I��0�]�x��w���T���R-�|�������s�V�0<�h+C��\u5}D�6�IMDL�C�61N����=/�?�/�_$庫���Z��dS��(�D�ʭ&�)%-����t�����j��p����A�|�r������R|{.*p0�kf���ܹs�0�- �<a?!�6[�2a��d0�|������{��) �N�J����V/���s�ب�`�=&�S+M_�(��6K��n>�t�W0�n
s|��-����$�	r�۝3Y�%�5c�N�劉B����/�$*������DSR�&0wp������j$H��@
Fq�'�#[�%�UK������/��EM7eRw'��� 6�-����~�B����n�v@�6�"w��<�w��(��#[6;M*��ЛQ~�W(h��_.n�I��|�]�ǽE�c3a)MF�9ٹU��?�a*�d'��~n�η"��4o���mŘ��5}��67MT+v�D�r���?�� (��U��΋	�k(��q��$��/[4����F�H�͚g]���`_(&(
��s"O&=r4+d��Tn�@��_�
|tS�\���a�]���7��54��b5T�9���c[�;�G%��U�E�D�A���g$���3�u��y9��[uԴy�(�,�[����qj�p�a	*#�#�Ƌ�Ʒ����(e��%�52o��;,`��vy/�Rr=�Ei��KUop��ǯl����m Yf�J���螔:D��|�kE7`�{N#T�H�zk�`�4͌�XĆ�K��~a�9[�/L��Z�\-�����(��t��db+�������� H�o�z}Bg/°�\�*�l���)k���v*~k ���\O����Ky�v�w��h�����r[�S��4Wt�I��y����r�7����*5s���?i<:3�:��g�ثYc����&V�9�{����ޝd�6# F[�Tb�"��74>c�rg�ea��!�V�x5��p�e�����h���d��5�X5�x�Q�)��r�{F#:!U�-b��xK>���Հ���{��f{3
��@�'(o�]�Z?�4g�����" ��*ߔ��9�
Wk��be=7j1����{64���6�|>7/2�{m�f�>~6^.�+f�b�m���/���s�e��p�]fǧ2�����k*@�ͦ~��D�c��`�Љ�A�<�F7�#��VQF�2��t��u���P��%�x�2�D�U��@�Ii1Ҝ�A��/�Ȁ_��X^3o�i�w�m�l'h�����j��w[;(�$bˏI*E/� 5��c�� �1�ф�6�`��>P�rK:0�2'ÅE1��'*�F������
G�藞hj�s�{A���Zk^?��v��LAy���O	Q���^�����{Ա6n�/Rj��(�i^��#�S�1`�u���Z�y<��]e2�L���\�DSR�X}T �_�7����B>�\z9���d���;^%���Q��v ��{h��4�b���o����:�-v)�հ^�J��X�w�9���.~U/��=swr��W~����̾�L����0>3�k<j���g�}wy��M�?#Bj�fi�C����k�6���f�X�h�d�.�og�B2H�Vl����x+�)u��\Pa=y��a.����"�{��^0A���d�ebgi��>~lڿ �w~�5bɢ�)U%��d۝y��^��]亽��IxԷ#����}᳧��Y�y�����۱�a8����uq���������)�����Ƹ��v��}�ze�:�4�&Q���ZX��?����c��b��:��Q�"�����N��R�M��u��2.�DU]�&�7��H��P'��>�qK��f$.ܣ5ֶ�gi���|�Ͻj�Uh�)F�R6��yd��i�����+�_�&)�D~F<�DT�x��G����[�W�kk���nF�=xh��_|X��shb{�
��TXV�X_{�7�Lx��{�Z����RiWw�K�6~Sw_�+�`h�����<�LJ�?�? ��%�:�aVC����@�k'7�����"~��~���Ok0���|~et�%���Ԋ ����M�߮�=�p�V��j���ٕ�ch������lom-GF��'���`yL'�)������f�K����مtb��
Bx�$���<�N�A��۝,�� #[�V3�d��	잧q,����5�v�tR�����G�J�A7s���2�Aq�3�H8::���\�m�)BA� Wv�[S��/ȃ��Ǩr��'�}(b��Es�B� � {��Ƹ~���@=I���8`W�|�(QBsJ�C~X"q0/|��F=My�H�������#:�b�����4R.�Y�{v`��Kv+#-�����|*��q�=*��������� �zc�����V������6��_M��F�5����v�;�{j�!W.t�g�R�t��� B�|Q8cj�R5�t>si��-�w������LJ�h^���k��=�z�9��E@��I�Ռhw�S�i���P�;u:��KDW��1����j��ꓗ�� �w�W�2��}	/R�6Q����o�#DI�,���r�sˑ<>���׌�:��!��Q����"}_ ��ޝ�PZf��ІV����ʕ�vl`���Z!��H�|�s�2�s2��@�s�:dO�o*��6gy���g��\5��2A�~����*0T��F���*���y�a3V~����T�.��ᣂ���G�˽�����4��𸡧2��8�64A�^��~y���z��қs�l���*�!E��a����N�d� #S�mf�@qt�����ۘ�X��Om&�A��I���Y��q�y	�|�*��_�p��;#���B S�&��p?�Ps2UG�yv��ѩ����&a��1p���K0 �P���GW*fZ��E��),M�پ<�R�/��V%��i-P��^S�]�]/=y�:�ބt��b�O��x���\��`����]@a�%��p��g�d��w}-���caF����� 긤,�6�E���08!)�h���/��0�q|��$��wV=9� -w����H˄�Í�\
���j�%��_1��cnDa�\�LpXD���{{�qrr�K	��r,����
���Q�d(�QE:Q���W���p�!�<y.n����R�K�+���A�]��y�.&�Kf�!�Wۯ����}s<�З<-�T{��x�\'U �sgy��H�����c�2>h=x�׋6�a.��U���슏���4��&�� #
;����x�q�36�3\1L��Ar�p}՚�R�iP�C��bo����w>��1	º��K�i��4#;i���$�:x� �';n�!���*�|'Q���[�y�)!�奋�+P�i�ٗZ�d.��T���Ɛ��I6V	{��=�ת8���$�e.��%k�,���?,��
8u����Uw�l���~��F=���`<L+�*բX< ��t��z�n�ɻI�� �5a]><,k�鶆g
�@\�$mz��h������HO��~('f���������G2T��6j�&}� �Kr�u��~��W\����m|I(�ԥ�x�6�zy�k�牟"�&�-����gU:���� /���{��s��퉬���H"@�P·��(� 	���s��V974�juqw'/��X��l*v�8s,�2<D��,Lk% �{�)�3"��	�j7q���P�֗|�
k$4W���]G�ߏXӁ�b*8L 4���5�����g��e|ʟ���N���=PB���,��e���|�x�Ʊ���	����d���R�C�mҔ�ql�	�-u���9F�c֙����#�I�H��Y�Փ�'�,>���SN(�{0�0e��Nr̡㐗�c�dɬ��-_oЩ'^7| -(������ {�t����
��L��Lր��g2��oGv{�����)��	_ Qg�n���ǴZ�ת#��wB�w՝��Z" w�e�Za���嶵�
��va��P �{' k���v��t��*D
�f	*�l��t�Q �zQؠ���?��^Z�Q	���ט���V �tE&���5\p
8��雌�4�G��z�FPK*��.!:������5Ϳ��X�����"/y���EG�j�YC�O� �o�zB '�~�n�>^(/J�{��Z2���IC[Ё��vX�੆�ʶ5����\�Eg�<�m����˕�2i`@A¸Uj;���K�/�)h��U��Z�Ͷ���/p����F���C��~3�t%	��gN�|F��`_��9.���k�)sPߝ���X�7���2nD�4E�d�߉��+�%7�X�w���C�K�~��͹����̫���#
�j�߬˸�+���� �ǮA:U�6\���a;��6�!��zS/��%-��#^ޥ8u��f��������|�4�Nej%k?��)�g�4�$vv�r�;��b�s�u�-D��Y��/Q*�G������,�򎑖�q�$9�S,Dz��d�Oa%hH|ǆ�xn�S>}/5���Y/|�B��1,�#d�QF��p�p�(��v�>_��F��ɏ �۳?[;�[�j���}��>�N)K!�L���Aq���Y��%AN��Ǔ��n�R�_��xU�kv�w�nK�
�"|�P,��C�[ �����1�Zm�r�k3�$K<�l�|��@�y������QV�T{�`�N�<$��ʐB{te6&�;��y۸���B���s) +sZdOq��6���@�*w��:��/3���Y�(���}=�$��+��ʻ?��bb$�[�sy�m�r�L�eL�r�}{hd�'�����IlީuNK�~?o1
�xG���F�Z�4��yO�|�$u�[��ނi���t�d2z�j9�{�Q��)��� �1�I�����L+��k��a��afb=�Q��nd��wc9l_Q�E�o?���
�S��֑q�οBY��.ף��<ҵ�b���Z0T���]|,�pF�%�Yl��{�^��.�ܖF����i:<"!�ŉ��e8��M�Ug����,�N��gZF;:��օ��+1�zm$���80\�k�$��~��B~N�ո�v���R��״�L�rIЛ;�V�<®ꔄh+y�^=ܗ��^���k���͙�;��w���l��Ls�Y�6<���o{���ZO$^���Oc[�:n�WCU�<����d�p�.P�J��*�g��O6��;G����~�}qB�Μ�T�m�*P��/�}ǟn�8Ud����+� ������+ �\�Yl�I|��߉�@�N'p`V�&$�f�<��A�'}�@{���y#���K5��C)��¨���9��N�YxT��Yk�	��M�*�L��E��%y�Wy�y瘿Fd�g:�1�����3�|b|��_?=�ڇ�{�BZ��H� Z,.�B�Tї���Jp���S�����R��c�;g�|�	�2����t{��W��7��O~���α��jQ&����LG if�y��2t������h�ž�t�e �+p��n�K`#��k�m��@&u�|P���Ωm�?��B
��Sj6�ULB1I��<Ҩj��-�;��_Օy�l-Ox��nݗ+��p��[���&V�k����-.�NB���L�_�8����=VdH�X�:J�1P���8��ˊFV��ſ�TU�-JK3�T�o5��+Q<1���B��%�w� 2�
���@���]s�!��^N?ҝ)��9a#��Ц򼙯ɞ����^�;���\�>�#�5Jnȸ<,�.���+�%��x�8q�a9�K�ۦ���&y���C����'h]k�K9��#WV��$�z>��`]d*���:��f��H�D,ܜ��O����:��ӑ?P]uhb�0���m)Lx>��}��UA��b@Ģ��Ų�*Px��z��	�8� �h�r� � U9�V���	ހ�Ye���� v";�^=�	����(2wG�eFQ��Q���DQ0�o�ϻB�E�ګ�K�A �_ŗ�<H=����9�9�e�S*']�� �ݨ���@�x=�]� Ǚ�ջ��b��d%f���T�#�X��f�p
�`��i#�J� ��*޾�Z#�=�t�����z�r_�
	�sy�P]p��g����ކX�+[�t����=�ƻw�?�$���dQ�:�[#�E@�x���nr�]T���*�ĉٰ�Y�c2�>p���8�D���-�2�'��w=�d�l�ɫ�<�����ȏ�H��p�6��}0>�+�t:/��J�M=�EXHr�J�h*� ������dW��:���cE���Ёi;L]?h�=)� ��:��t�M"\"rGĕ�>�>,�2>�����+r�w�n�Z4�Ѯ����W]~F�Hd������kiq����<�S������c�hi�����<ٴ��$0���)	��w��?��3�؎΋E�`>+���BX�("��N�R��(� 0~�z�Ä�{�����x���w��C�Wl�9�fQ�&2�� B�l��z��/B�}��ŏH�W�Q�\�W��UQ�@ ��$,(��=H}��Ɔd2�p"�T��4^6��=U@�d�?���.�~{�8�+S̴^~����YI�W��3�6���Ds�.�~�~�����y&�+gY��J`�#K�^	i�0����F����74��n~P�h~]%�����@\4wH�߉��c�S�Z�*�L.--4ZS��V���v�1Q�K?P�_F�4N79!�M(����b:y"�2e���;��(Y���̩O��=�.�^�
���ĵ9Y[V�
�ԇƂo:�<ғ5[��>�����y*RH�ե���[;e��`�n���T)�@�o��N� �)�ͫ���m�Vbb�{g����ྖ�.csD<�R�{�h�ʂ��X7��}5Ho��j�`AR7m�2>���	`c��`z��p�>��IN����$fy��C-�n�^���&�ː��Y���z,�Jf_`o�R`�������Q����V��PYS��V�Q3�h��O��g}�����e �y�t~Ww\R�Pwf�������_�"�Q�6ũ>�Z�������o���r��~ݻR0,�A�|T�����3!�Q�['d~Ą�v'y��!"f(��~���[>'�P��L��c�#'�AP�3�P\?�t�X鬇\�v0Paw/�}�odu��^��KpC��W��%?����\��f~�xY�
8}wz����;�������"�E�'L%y�DӤ@�q�U�3^�Ie���L���u�~]��dF'Jჩ��(!&�u�p�#�}{_JrВS/ۄ���-O�z��W���
���3�|�����T�wd⑸�U�i��ؤ4嶒���,��f���vN�7�8����������fמ/ �O��p"�?��$%���e�f4fWsA��R����XI�l/\�(�B*��Ε`}0�������I;JS��з��}�v�y9�i�f�Gӌ��5����{��z}��� �7�fh��T��A�K���zubΌ�7<&�4���	�h!$��Ŭ1�<�a�	Z��»o��W�����4��m�V����uFE��yzS���n�Pj�0i�HS���N��2���.���s������*����Px�I �35���wtN����<f@�n]�9���e鞟����c��Qr�I_��U'{ص���� �mn?���쾚�����D���9����G}Qz9��}ó. ���];o�<!9a4�ع�]��gl⮗�`{M1�R��"k�Z�2~	�}Q��f.		���Nr�aߘ:IS0�\ _vo�������&qD�{��(�Ч}l҆_ B�ܦ���tbTK��FY�"�e�(��l���(`�ƃ��JI�P��=�1
��5i����t�pz�d��'c]�_������I�ZZ��o����n+zFۂl�Wp^�u��W�*�A��6����(��l �Kw��.:�U��k~f���? ��ߡ
���@���ޣ�xRfz���9	���V�bL|�1�i}O�s;˶qp��O�������Č/S@���BO���:���a�}�������-w�1/��1�X�-!ކ���)U����{}�zP���T+K��x��̜v,����_8;]:o<�^D
h,���Bg�����G�u�ۙ���T 
�%x�A3��ǂ	��%��	��^.����	N?~S$�Q֧�V�1\��D������v}���
�����|�*w�45�T:��YъG&G�3�_�̤Bl��?D{TC�Z�� R53=a���coū*��?�"M	����.S�i>G���vSt����z�@�G��n�J�n/�i��H(�\b�$o�E��d�o�?�G"�h��&^�_�Ў�m��˹{�y��W �Y�����p���}�鲳���6c�+ZHj��Uv�zF�3�����Sm0|�'$�E�����=�*�f�|�-��7a��v�%����o;�j�A,}�Hd`K7�M������~���(��O6|��I�z��W~�R̶v49�e?�լቑ!O)���Q,+��ϕ,	�n+?�^��B�;UÂ�n*vڈ�M�h�"O4I+?�p��)iLc�P�R�6��Z�0��d�]�xP���"��T�ר�*
�{[7��0�5N+��V���$~��Q���:C)N�}4I$61�p�Lr^\⫇+��ᯍ�����ǯm}�6�~ۢ��u�	�onі����|} 8��~���[���.�#��?��[�#�L�ɮ>��E���)(�!��x���Z �X>n$��7ѐ��
�ru^�\k����{7�!�)��25��x4Y	���y%*����������eHU�����Mr������:�[��3ԍ�am����fΔ�Gh=�s��ӹU<S�]����ɣ�Т	�AX� �m�lm}��q'>��$��.O2�^Q�mX��=��7�ݪ�-1�ͺ�
��ȸu�&^��Vz ���B�z�������0��y�{�*��v"�ܖbD3�$��K���9�tAӀwM���,WAv0~��D'|P&�=��,�n[��hչ)�ˑ�C
� ��o~niρ��dv� +<��KT�.CjC�����a��i���8A�MϮv69����M=�@?�W��3-���%
@q擏��Pp��w��׃����1�[3=�%˘���n�XM�78#Q�e3.n�L�8�Ј�2G��썚1?�~�O� (2x1��| t�Ћ� ��,
^~1�a�*�0=!~(F���=�`nxK&�9�H�[k�j�<y��S�r�{�y�B����v��i��}��Ǳ���ms�O�Ƞ��R�Hk���ލ䫄��}����e��ní�u��4z����`��P��0űxԵ�O&�����2 � m]�=�T�D)���s�T�����[R��kF��jH%4iI8�@43S���!)��9�����Y���r��[�l��2�\^SPrtA�yB^��x�*H�P��r�����MO��o6���{���)+�J�W����}��R;��K��/���٫[d��s��t������ާ�p�ϮAk�_�g$M�����J�EE�%�\�4�7E��hQ8�M��Z�=&�j�0�V��5��"\J���U�|�1�  ���g�0�8Y�&�;,R�I����;���^K��sK�._�;H����c�k��'�U��5w7�DH��q2�`�UU�	Ѹm��n[�K,&��� �[~��sI�h�R1�),�0��q�5�<�v�x�	Q/
�:%������%���S5�����7}s�k"B"a2Lal��᎓z��f
���/6Z��;�DVġ�}���+C]�3zkr!KF�S��8x�ʕ/�a��S��X2y��{O���Mg��7���:!]/)S�?y��|��a��;�f������B�piԘO�,�zz�����gY�c�$�ze5�;)`���-�FA�R���
g�V�6�-���b�(�OT���ۅ��vh���z�Aq�;���m���O�Y�̠��<nv�$�a�����1�8�FD�Bc$P��ke�t�`'ܺ��oF^TT����:k5��y��K�8(��rV��b�>h��Ś�-�h�\�OC�z���c�᯷���f [7^��3���m������)��+���4�|Q̚�π�c�F�G�k�y��'l�ϵg�q
��q��񠲲�K!y�֬BH�bjԑ�7�/�Q_s#�6�	�F�vɩVx��Vf�kM�0��(� ),�s�^o�/f��򒻋H`��!�bqe+���\�)�{������+MR!�qx2���A�6�Q�Ui�m�Np������F�B�(8�y]����%9�
�����f'UBѢ�K���0��Dc]o����~�->�M����<�W���?n�	���`D_��LA=6���èx��EX���tR
�L�����r��A�N���������d��\
�ܺ�7�wף�8���G��%:ңW���E��#������#���=i�{��i��֘RT��	�m���c$t�9��q����2�9��#�	��ue��G��τe�?Q�tf.Ψ�N��r���Z����Z��?T\ه����od���9��:��������7�VݔzmRm�UxH��;
#�� ��H�|XH�������*�n5R)t�c]�V�̾��M��݁�P#t��=������X�Bfh<��D�w9�p���6��ʥ��n�97���h�^+�ߜ����3�ϸ{t��#�Z�@x�&�Czܽ��`���/kgI`��}8I_:��A͗���`O��W�	�Uw"W>!i����A�Z����}�ؗ�&`@u�x��*��E��c��,&����4a�����tx�i	L�=sb�@%��_s��y2N���r}�C|a�SӀ��|>�Ȯ�U��.j�xJkᔣ��p;й�D��J�P# ћ���Z�؞��ϢR���ZQ�<E���=jY`�@�	=�D��=O�=`,��e+�R�I�D��	�d�T���ݧq1�e]eCnH��$KsI�����ʒ�w�(1rӣ\�=�$������ݔ+I��Jd��a\Mۯ��;A@k)����&5fU-˪�w��<&b4�U��y����P����i����j�ǋ����ِ~?�Z5j�p�᧧�-X,���`�l�ΐ���&�QYx<�2�I8�d~Ր%E\g�J��=d2���&3?qj��;y��#�m�ik1"o����U����f�=v��	��ŋ*��y�7�>d���NY��3�׮�e�H�F�
_�es��=X��.��D^����U�̧��(�7���Tp�E�Pl��'�0�hDZ.�"�)m��u�X�Q�����x����s�qƲ~�}d�f�+�A��ۍH~f�~'܄M���}A܉�rܕSW�9�m7��ò�8���dQ֔���s=G��V(M]�����=r�w%1�(����"R����Wl����h�pO��<0V��un���1;�W��s�f-IJ���+�����2[A�����@���}�����9�`M{�[��۲0��8�'�wS�o�y�=_R�'�@f��C"����*���S?ǵ���7@��[{?��n~! 
��$_���R��>U=,hN-��C�n�anH:�0���^+�-b�����Nſ��:L�G5�e{�P�� z� ?��-�NA��X#<>ݸ���۬3�������h2Fب��|�[Mm�k?�.�\����xk8�H�Q���HSÛ�
BMЌ�p��,�F��Bxl��Zt��i4��w���=�j��լT���	�F��Hxx���6	4�Ze�׹L[)u>��h�]3y��O�m���k�*��z�`��yz��q�^�d�v�����Q��;�$mr-�
 ��w�C;4��ݾV,��bS� ;������#DI�2JV%A7��*Ҙ����ۢ�8+zǇ\UY�!x���8�L;��ͯ��҂��_G�Z:\#�ES
In��]�R$ä��5�i0Ǖ�����@eW���T�U[���^XkS�(���l���s�Y���ϾR&}����|�M�?�F���a�/�'^b��)8�c�{��*#`�L��^��v���'=E�L�ۅMcpԜY �J�+mEr���(ӝ��]�2X|��`���F�����U�YKlh�oBuÍ孑�B�ߘ�q>�2XȖ��O�P[������Z;�������&Eh�#B�7�9IR}���ɇ-	���� �n��+�r��1�n�#�M���\��B��@�7U�O�͉fb��[�+X�?���V���69�H�|Ll����S����oصv��
����=ԧz
��E�d�i�=5�Y��Z��ȟ�M�9�Y�>>�{q�1�#8u��`���9�a*F���Q%k�V��ZJ�%7!C�"�,o�_*�]��Hя^����{����w;��Yv�sb�^5��K��*h:�\k�P���aVF'��%H����^!����l^`�����W�u��(P��Y����9ƃ-�_0�C7�ؓC���ڠ0��A����ƀMٍ��W�r���[��s���v��G�ߠ	sw*��	^[}�B�����,^�x�<��rԅ�F�l�0GXF`��"�l�ڊ���a	�~lL�j�q�p�뱑�� Q����#�X衡5� tRu��+�����r<wj�X#x����M�����I&�:�a���]��!=U�9�,6�x���`�6D�QvaUͬ�h�$I���Z{�X-�]�A-♐�Mh�C=M*+�#U��N���}U��f�c�^���	W�6��E$��Z l�ds~om�v��Pb�]�d&�'�	�^ȱ�+(��5 ��"_�q�Ƹ���n�x���L�RTA�;��I�O�7B�F��)�]*L٪�v��W+%۬��Rs�-}�|��:� ?YV�<G�1����ޖۢc�b�2j����'N�܃g�:z��;!ՙ�wG��(!��8TgH�<m�~T�����`�&j�rk["��ł��6@�a�#�Y@C-���׭��i~�
��Ȣ#Ѯ�XG��/n���3�S]��cY��=(���7������\��Q�U��<nշ�R�̣(�6@ax�R1c���0�������_0�À�V$�BRei���`<�%]R'д�Y���-�A�*�B��"�I���P���\�6�- ��V ��?^~yC�o*I����Φ̙��s�"o���Dh��Cd�#���)/�j#m�r��0с��b�Dg=�Y��'N�+�VM���h�ȼ��.�\�E���k'X�)��<��N���0�Hy`9GN|qFQ���� ��t�1�,u��'%�ɵ��O�W 6G�CGu����+�E��s�dȡ�f�L%�F8W���-F!��g�����_6'��������}�E�O��`OkӘ��*� �k�mL�f��%%��/a�6j{�m���<�c�����?&���\����j0?.N�B�E�J0�G2�^i��:/]a�s�E^�Z!&�]~'=@P�����6�A��t/�0�E�!�*	�50�Qƃ�@�Ȏ���ӗ�H�"����פ/�B-��ؓ
5��!}�5gl)�a�J>�,^j�Ch��Suvi����a��Z�TYR��:�K%���� :oU�L�����F»m��΀WJ�!H5I+�`�O.�س����0��5=ha��^��4�kTS�x=�������.f4M��~�����x�3E���.a���&.�`9l�x�V�(Q�p6��G���RQu���"ZbP�c��Yء�΀A�0Pf���ؾi�ʃ�p��-(�e�� |m��'����Vfk'	�t^@���r�at,�_��4�r��$~<�~��{�aZ7LD������E�.Ƣ=�"�YA^=�g*�a]����3����5���$��G���bϿIȯ_���AE��i��x�D��
�Ƕ�i����V%��� �M2����+�+f�wa-�a�xE��"���Zl=x�Xn�婪Sp��Ptq\<��-uA�p�G3b����@fww�S���(��q�+�\Fo�7�&O.��t�
����|scFr�ôl�4dJ��ؼ�m���\�L �_��KJK���u��%	�OTڃ���o�i<�׾d��ڡ��GR6����*��[�N��u����9��ƗE�]�B�ؠ�⚨4hm`A���ި�s�w_MvBr�b�Cл����w������f��wv�9�����^�#�icq�)I�p{��h1p%�7���t�����
L2t
���$/|L@���9tJ �������<�$%�Q����3f��˞n.QW�i����!�����B�񙆀�O� ��r�(Q�A�C�k~�D�GUh�/ˆ4�w��;[�t*_m�s{4l(zFr�j���}���<8`ov�Գ9Hc��l����CBQy�>]�y��vBҘ_<�k�@�v�?��͖j�"�{9�#���.�Ӂ-So0�T�b
���*ћ�$ತ֋���qU�.pN�Q��`�q$�T� i�^���g�>�r#��>�|9Azq��Ͽ#Fw�6�_�M2��}UMc($I��6�.H�Ĥ�v?�T��WKz�L��z�ꆯm�"�z�}�ja���<�KV/㭀���]�b ��t�� ���Κ�=��/��j؞ϧ I�bd��<R��=~y�v��\�S�\���j�2Sǧ�������jY�)Y�����t7�:
^N^��4W�o{��.�Uj���7*�	6Dr䱨h��=��[Zƀ��<n�|?HRG����`!�={�p����?)��݅��V�}2�oͲm��y���LPE�u �ߝ� ��g��<l��F_���VM	TK<�U��`�h�����4����b�b�_^�5 8	����s)��3�2�6����
�ZS#�t����w�\���b�SF��91`����e�.'�9M�����{�1�v<��r(S�K^(�PP��9�T��{�U�P~��b�!�@5Gؙ��Ф��,\�L|N���H�,cnq`0�~|�sR�������g���(�}��:��-u[t.�M�.7���x��ND3���Ҧ��`a�2O���u��FCH��s����9֒1%�8�ޑi\tT~�V�*��+y���]Az��IY}�Y>�^�����ڴP��&ޮ7n!]��w��[��D1��A;5�o�Sv��*��{�k�䡶g�O�D��5y��<���'�d	�����]ŗ�|� ��z�,n�.���;�8�K�)���G��e����F%�@x2E�/�ަ ����X7�!J� �">TI��*7����b����i��.�p�	�V�I�+pD�Ϗ��!�V���2�q?[%X��}�l*��i��Jy�<8���}ih�89g�*ux������ �o��c���>K⋤o(l&R
~�br����6�'N�#��*�����1z�}|�����~�ՋT�u�b��X�ޤm�q�ռ�����X���2iDr��4U�����/�R4�Ł�cv?G�.Ps;�d��#�]�ɑ�v�pc �[`lZF�����08�V:����9�q�O����> �0Q#K�̀�N��Iഁ(G��b�F�ꤗ��B)���G�q#"�TG��0���:g\�іѴ�Y�׏�R� !�\���Hp8�ŝ��_�>��9�EA��Sc��?�47�����ה�vf�G���&H��e�'^z(a���'@�0=ܰ55�����f���2��5���Z5�;W��ŮJ���s+_!G�%d�d�d���"�Ѹ|���9��2������E���æ������d��%��M1\(/+��6���%��H��0}��V�e5��	/��G��2�rP}�������?N	�hV�|M�:'o�?]�l�m����kC޸z�ͳ��4ݦ oC��I��q���п�!1�J@^Y�.�oVf��o@�dڻ�m6��]?P����[��s�x����e`�B~��I��V���3N��r�o��=h=�x��'�#z @�Sm��gN�oX�����+�U>O2�ƔMB�n���KaC�b�~L�x;\�~⡲%��ߛ?ks�V߮E�7i:a�(#����7��<�cn,@�Q�R���W�SH�F

k�Ġ�)�j�?[�ޠ���j6�0��frb:V���w9Z�!�[�A�_5i�M���[V�|��Ӎ8�^�����$:�$8��jk��:~��3�_H�c�uu�I�k`�.�б_�k��Ƶ;�z�>��壙S����Ggw@U[�7F~qY0�!/��;x�K>#^B%h_:��Q��8��%Zi\Y5�鶒�9���4ˡ%f�+yjH�&����"������a�Ձ��yi�r��p%�)�Y�k�..Z�Н�Z����8|	-qIS�%��-=�,s���cO��m��9}��>��/3=ꩰ/X	k�#���P6�wkv����}+�8S�`K�(��H�N���`F*p��
��N�]��wEcΊJ�Q�j�H ^/Ѭ8�����>%�5���d] c��-�'4�6Ő��0}� �����U�xx{��b�ȯ)� �^��`}�7�ZC���R�&��*^M�C�5E'�d=�Rri1.���O������\�a-�^�F�������L���r�-�I�c��Ix�_|̙���.Ũ���Q�H�+��3�� �<�9�q���k�P��Ӗ�e���f79Y�!~n~7�E	��{rX�xk:����ѣl��T_B��	AL�0$jN�5�v�8��*%��@h�8�u��X[��B�$1�y��f�؂˜���E���򯱄^� Lͬ�r)�I���]�%�N��7�[��v�<�����B�i-�D���4��* 5 �8��3�pɶC�SA�_-�q��?ix��G�
�ϘZ�Ե@P!�f�u��>B(g�QJL�a~m�j{���zL'GMe}�,��[���B��y��aZ(�i��'#|��h��,펹~բ.|���
�4��	�2bg�^�j;̈́G>�G�{��Ӹr��%�i��m<a���,��y��&�ˁ��q�JФ~b7V�"�)��9??mm�2yt/X�z�]��өr��R��Kg6M�5�O-�M��[N�����q6և��ss�~IO�u	��}���X�zzDZ��6���x��I�<,tԾKO*�w�<21OP�v͑;�*1X_W��֎G�9�9�[`��)�Z�Jy&X�լwj٭�Ѓ-p��y��|Q�����E������0�w�Ȗ^��o{���+� �ֳ�mF+`�֍�va'K��c" ~s�8�?]_�`(�^X�I���p�A���2��3]RIv�^��N|G	Ԩ��o�e��?�&p2�
J�X|���<[.���|��ӥ������p��_��2�ɹ��"q_�E�ց��?�X�r�Jp�X|v
:��X>{��?hQ{��+���I�Vu٦��=���g�(v�wXڍ@��l���fM�j��&�"��跕\#�gB}š#p��Ng�oC�s�t�:J)#(9��+\�$o��ɢ���6'-�Az���O�0�� ��IJ�����b���%[-U}
 �`6���� ��c>t�ó8��b��pޕ��QÍ��q;Ru;l�8~�~���!��S�<�����jW��]&[��=*F@�%g�N��<����fg]x��S#	�$
���w#5G:�~w3��|�+yb8tK>��z��"XM^^{�4v*^�A���M�H�=�@�7��A�ę�G+�W���~> �D�| Q�6a�Zt�Ԛ�@Y�\U]^b�pvݠ2��< �0aq7һ̻�����~L�߽�w���H�`.���������F�֜�J�h�akS���=c2#7��~A�_k�jir�+U4�7�!��6����š��D��_���A���:��fV7�&���dg�n}H�h8�L �ͣ�q*%$�������[mq�`���/�����Cn-��I�!9��a@��,գ/o��"R��z�w�-x�]�s *e�!��Q�ߍ\�T"zd�)u���J��0/Cn����<��<�A҇?{z��r���5��Ȇ���S�l�Q������U4r�,`Ȣ�]�'�eH#�lɅӢ����
��M|Vt�$�����iD`�������
c�\��lּ�D�yC���mn��#���c���Dk�C�ڐ�; �����~�8&�`U�~+��Q���ӽV�@������8A1yݦ�����I�����X�q���Ƭb�)�<�&I��Q[�<%&rɹ��ˠ0aD����c��J�b=m���U�{3�Tn�p�Qs��%PNj��7��G#rH'+�`��� 55�T
��/+�tW��4h]�<߲�z���O��AcъPpj�}M�_�{pa��5��iZ�n�iI�A�ó�ء����*!#x�zb�b�<�J��E���'�#�'z��lUv4�rVn�X��O�g�@��ވR����V�FS��m�^�U_dr̡�"G�>�����fp�����M
DO k��q�FD'@=}�`<�p���`��_GV����8�K��P����{�H ��@�������?4��/��mV6-��G�9���+��0�R\F]�EaD�sv�&�D�pٰzӛ�D��@�0��"�v�&�o���%�(%�r:;��Lu�I�Ol;�B��'�N��������ŶiJ<�\����G�K��Vq����z;�͝8�����2&�uе=�}.�ZB�%�@=�B�����_������u~�	GLw]��a37ú�2[k/���#��#�í�n�m��ϝ�+�g,x�����ƠW��6BO�V6a��\�z�-��Rbn�������UvR������&��x�cZT��*�.��[|����WD��~���\�Dnx���:����y{���h����.�`Ij[$_w�ir�խ���_����:�&BDy��٦6���ک+E6�� ,�I[���v�䰵j�A��^��%{W�2DY�8*��I�M�����]^Lɞ	`Y��f��eO�ꎂ�R�ԥϛ7�6����U�5�e�)�]�9o6I=,�:1
�>�E2��Vm �38�?��\�:Z�YQ���������D�U�z��Gx�7����s��-�I�v�bѮ��dx���V����c�š��k�t�t���n���"��Kp�Ȫ�r�O�ae�
������1JΈ�=�!���O4��=�?�n��h͝B�"K���`���ܮ�>�D'������Ip�1a����+t��|X�ފQ���%�����C\CFK�~sw���2���@$�D[���y�/��=ڄ���Y"+�5�7v�ß"7���H	��i�#��^�"��5���������H�ln���'5�eBg*b� l�PC,8Dp(~��@�i[Ƥk�K�0��sw��:�����=����y�����C&�CI���~�Yx7!� �Ȗ��<� �Mp�?n]����g�/����n&�Yu�N}�S�Z�˚�w)���y²�N��X��{�-?||t��	+�x��xn}��>5�Ϭ�Q?��������>��D��yFM���VE��}�;�'X3;�