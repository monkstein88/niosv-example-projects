��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a�����/�	v�+����@ɧ-3�����Iz�t�܀Le'H>	6"�U{��9�bEɤ6-�!�V��s� ���m�|����~μn���}�iԹ*VC�4���m7���-� �7�o�d�0w1 �⹺�)=k�:+5:� _M�e�$�"��O��0U̅�iZ��x�K�~̏*���;��R+X�="+$Y~�ml���n�H���K1,���0�ϔ���憲e'oN��D_lxY��^PZ�#�C�e��Au�֝��2ɤZ2���ܵ� �o���ǣߜM0ځr5r`D.ɩ�
e���
�Dc�����gC�8$����lc'�'@��A��Se��J�oY�\�?f�ᕭ�o0�\�O��H�$���m���M2�M��J��?�c��ˈA���~=ɮ�����D���B�p��;�e㹽yU4-����_8����p�R�C7�H��;v��F��5	��zMV�I�xB�cȀ�j��� l�{�I�e>;�IT�NF.v2���hb�]%fzy�0���#�%�GNאsXU�թ���*��j�5x
�P2V�?��9}��=�->���x�/#v��_�����J�N�(��x�USy��i7�4��J�ÞQb���u����V��i/��R�	J�,W��r����tx�E�r}ӣ��בrl��P=��������1+�&r�W]�#'`��5]h�?�G�i��:b�P�Ǎ�;�׈6����r�R�����
m;��V�j�w��^Q�Z1�d�p#��`�h� ����Ҹ"���'�1��o�}��d_��0�^$-9S������b�I'Ѿ(==� �����N^X39޻f�z�M߶�>m�84�G�d�|6� >��2'[�a[g� �oL�(Y�h/G���ܚ�ղy)a���l��� �d�,�f5�gFS4|�M8l> �����0<O`q�`�U�X�$.?@�S�xm���h*#���_��)��a��i��<g��Mە�����3xt�F�����ef̌�����:Pn�� EM�é�=����/�̣S1��$��<a��\u�!/�\����փ ���:�u���־��Q��2�sƴF�X�������)|=ZϠI�2É3�K�%3ń��q�؍o* t"it`�+��7��܌�G\{�ף�O���Y���� �i}�{]�u/�{��"���>OL����: ��j�3?/�̭4�c�-:���;x��_�ѽ
e�mN&;=b�Ve�tE�;��n�1������I
eU� Fo�#
I"���j����J�k�jt�G�]3��у�'A����|_��sZ=j�֔��57��X����[��	Y'�P����&ѱ�iQ	7
i��F<�|��|���i�c�k@ߦ~����ȓ7�moy�D��佻?j�����**��ڞe��ܟ��1�DyF��@Tz'��H�.Ea�׮!�y�ٽ�!���FQ\�Χ��=���
Vwu�q�s \p��Kȩ��>
Ҭ2b����9�h������'�Q�}�\h5�f�3�d�\,���\���y��t��ÿ�#�Ⱦ��v���^��-�m;M�:�S�P(t�_e���<����_O֜���:�Q
U�(5��QI\��%\wg�h�RU}w�^�sT2Ĕ!��WDŲ���x����f�'�3>`�fQ{}��嘝w�;�6�mo��Z�x��U"��"����;/�u��L�=P0�4��#�pˡ�������n�7f�����U�#�DD��<K�:���&h���~���F���d��Oّ�����v��k�Kō�5HU�@���`@uеh�.2�{A9�'j)��^Rc�	b�1�{���~��.臅� �g8@�"x�_�W�;�w?��� N�O<�>�W1#+���yIyFCBW^ج}��&�l.?��}��9	���Q%�8'�(;���jn�0�vp���>���(*ԡ�A4�WGr���Y�w5��+���bCX�N�<���7\��b��)ee
L��h�����'neĎT�	$�P�h��O�� �n�ު�P�>j�h0em3��c����<��W�pT�S�3zН�eN䎮���1:#@&�*��K���"�_���@��t�M^T}��\�)^9�W!>f;�Hr��}fvx�L�:Us�7f�:����*�6��ȩv�-��X%�F ^fy�:$�vr�n�*�]���^d��3d�æ��2�1d�.����Ӆ�Bg�H���x9����ۥ�u�y�*�*��stc�� ���*V��w��쇻כE�@]$!"�� ����n�	I����ľ���X�uZ,�C���E^��S�;�K�?�X353,��w�����n��K�����x�{�
�mu]w���:_%0[��YOIgp}�ԑ�fh��w�nK��@���=��V�V�fQPD�8h>��lx�N�8M2��� ��{ͦ^��4Z���N���	�G1�I���&̑zU�b�ޤEWѵ;���km�Г��.���]��oi����r�7R��ƙ���b��:�.R$]��M�(,��T�E~����t�u�[!X��ϧ˟�S���rO?W/~���|=
UC̅�U0���rsӆ��I~�����L�f���8,���0���ʩ����*2��ﭜ�h�#3����$qew)�aEGs��j ��=��93QE�\=ǘ�P���X	P)s�Fjm�0o��f����Dd���&X��,�־A��p'0h3_�dc������]�FWR6Ҷi��՞��g��$z���	P�q�mH���k5$:�:�zW�JL�t�3tg�S�Cs҄Hg��7�l��I���ĝg�4�\&���l��{|�uh/�V*�W������ֆ)���Ks/�)Q���-�q�2�)("���D���1/L�GӁqC�#kK7֜��=�>\`��ߵC`~`Eb�YvMӫ>
�hre
�%�#}�of��r���/ �'Q���h��/�6��*�:3Ǿr�ڑ����[���pP-ӊ0�W����5:q?H,�q�r��}�Y��^$K����l �Ӆ�`E>5C9o�ԇ�JjE�{��0�_8N����ZW'�jQ� ��8��-�~�W]�ׁ�Z@
��,rt%�jp �68�W�X��&ɦ�8Lq�=6Z� �s�������u迻 Cy����<Y{�.ZHxJi%윰�P�)��[E����۹���D��V�m�˶\�t�4� �Vۓ�U�#juԀ�C�H����1o�g���*��s��?���p��u,�+,FV{�z3�Wd�2��>2���3y�Ю2��[~d��abS1qn�lq�^Y���g��=���e���|*4�7�
~���4�D��h�D���I��#�[<����ilp��NԽ��R8�#�r��5���~�
�%ޗI��ɜ����
lU�@�U?X5���ط"�Q���ER�jX�+���K����9��y��`�n���h���p�Z[�iދ�˔/S����]��kQ8Q�q�U����[�@�RA�c ���O�PduZ&���$�7�x�G[�j�.��׹y�r��Ɩ
�{�H����ͮ�t��>�g�D�I\5�P�p��;%eз�*���26Q,�"-܉�����Ij����^�1�V[S|\Q���jA��3�C:
%>T�ܪ�Q7T�4�c&���ѽ���G?e�91r�f���lB { �s�L"�E�x�;g�#������%s������W&蝰���������z�:��sڽ  э������̀m�V�S��s��6���M��b���(�j�_T�i�k�@��o�!��Ҧß�=%'��+6�W���@@0}�~Nɾ��5�a���a�h�݈P*���{@/U�!�¿� �\v��PMΈ��Gް�z���fo��ʋ�01\�5�Q=�w��W�zj�	��-?11���̈LW8�kyV&�b�[�Y�&^�s�B<�M��p�>�Uh�����sz����x��K9�R/Q"�r��֝��O�UB��.�7���p�)�q�g���?�=���q�`�.�М���Tpw�Z��[y"���L.;+kë�ƫ2�m�m��Z���Ѩ��&���y��ƴ�� :��2ҡ��� �)���ॕO�{!m_ϒ��D�P��2�� �Ԯ( \�\�w��y
,tV��C��7�<^X#jh����S�Lw��^k~�7���&{!U ��XH�]G�;��0���B#}SS$І/c�T1���UE��g�6��/������񪊥Q}�W��Yd�9�&��P��'!9`t��ҧ"L���᰸�F�p]1҄U��!�Ip���af�H�H�8���E�qs<?�"��RA :�����t�/d����ِ�j[٩{�K�$x7�Q�J.b-�+��x+COE��L���.8�<����`�Oր �(�e�;��ALӍL�?��h`h�F�Ø<��Ӝ婆��W��c�Q��SX줯��K��{�C�Q���|����: q�Ģ���Z�, ��0��0�.�X���ѽ�9A.�WA��f�&�q٪��F;B��З�@�Q3PWI��,��U���P�R6���[SV��_64ޑ�j�*�����ޒy(W��W�:\ZON��D�E����ʜ���y��ᚐ�Lou䇅�mb�2Ė�G�yrj.�}ܧ���Z �чh�ရ��7s���k��� 5��Ѡ�)���i
���a�lZnd὚�G�~��ΞN����T����e��犫���xW�`,֤E$��*�9S��T�����q�w�O���E�4�������I�Ȅ%���ȱ=�\Cm�?�_���+���O��v���x� 2�M�9��&�G��zvL�5
t(�����������A֝��Qx��X}9�7�Z�?��NCa�u԰>><o�3@9
v\2�*�%$��%5��A�t��������v%-IK�	V�ܭo�+nל\Fkbz���ӹ��I��|��1����ز��5ؙK�~>����teTc܎R��c��ϑ�.D�#��$~9۴T��-�/$XuF��]�U�W�a['e2���-^$ٯ�	G�����(�u0 ��/�;�m��+03�0;�"*��
��ۦ��^W({Y={�G���_`ӜA+"26|l�U_qS+r#�|�(�Z��T��/gv�[��M�EL�pA�
Ѣy\��Ԭ��P��!�J8���<P^�-�>"m�z�35���$d>�A����9ʕ��q/��5y����,k��>��t>�s�C0ň��Ȭ}!�
/=�#X.�V��H QUl���}�����c`z�9x����X;	��~���Z��i�bHPQf!��[e����3^���H�6�+p�V���'1*gh�ʶma :��Ҝ�/e�Y�����,t��K�O�'�|�}*F}���R�W��(���^O�$u#Ʌ���"���=W�T9"S���#��O\���"@������p���Ò})�P�.?%���hH��F����$�7i���1y\S��k}'u�h
B:vM���&�1_(�a�Н������{����U�"�� W��3�N:\�: ��[����z��o�S^8`p��e���'�
��Xa�}�PX����;-#���TM;ץ�"a���[&�z1ڋX������=���<�H��?�r�_��dMQ��:���I��v7��dm�_KX" �c�������=�<0O��C��t�x"+Ba3��D'��)]1�_j����k8c�S��WP'����}�:�R��}
N�}C.��c�B�k�C����}�X�]���ՠ�ʊ�)�!�E�c*9L��o!ts��j,y�m3}}U����Mǘ�3x��
"X������
�|�S.����p���w�I�'hv�yH�83�{h��BE]Θ��6��nP�c�	���V��U�7�A�3A[�.R��3���Q�ɜ݄��o~Ր\'�����F��I��4�A2��8(�oHR�- �F���ң�-�qc�;��E=3-��ǘ�B?vA��u�<0�`��(�|�m�VE4#\<�yK5#�[H�_m ;1����=���"P�5����BɈJHP�z����Uc-�>�-+$����}��.�.��4���7���1��,��XA���	1��z� �>ku!:8'�&u�tV�v~Û��{�=���{J�"�Q����ynAg���p�p�{>�_W�H���4�$�ֱ�$s��g�x{�%��X�QlR���;�1+@)�z�o�[���G�Z<�1|���`��ި϶��n�),<�^�wu����F⾶�T+c���[�}g#�~��:�̆��@h�Ҏ��3a��c��~���b�a)��l�ët����(��x�N���8w�H[�KM����u�'
dՁ�=�(sbpgj�Q����5�M[؂���\1�>�`�_��aR�?ǐ{�7��,Fr�:AXW��Ah��F��;����I�6�<O��b�U&�l}wa&�>&k�rJ����Zl�Έ�LdIF5���p]s���mW�B�� \��G?�{�C�[����ǿ"�٨����	i�wG�tx��4u�%���\S�	7V߇>�d��DȪ��-v��|�dL���hi���l��_[>��[�sa$�Z�jcя�)�;KW������� ��[��ˀx��*��/1���L��:H�y7-2�-*3	m
�P���݇$b�#H���:`�#ň0���D2#|����w���'LXŏ)a�Z���x �p��?{��9�5_���+����t�q�zm7�K2+q_�'7\\~`FiֵT]���높��n�6�Ta}��/�r\,6�R�W?�l� �cY k���k�kz��/#�
&m��A�Aг%�5Plci���>t�$f�A�[�T���)���vκ"Z1(��i��0����io&��N|�`2��#�v@�'��)ɺ_H�/�/�uՈB?��d�U
�������MT选�Ѕ��#y��S��)(�ɺ�������7�C� �h셱!�:~���)\Σ�O�K%Z��أ#�����D��9�%�T�:��<���׃�5�ˊS�����i͒%T6��6m�-�S��-��_�Il[DFq���{Ud��S�@?�l�{��Mġ�[�����(kk�����LJ+y�#�5���oM�܇��Nyڦ��!�+l�X)'��İm���^~ �L�sV�?��ni�z�t�����dcC��.��$��/����Į4�K�I��nZ���SW�ǡ�;��Ҳ���3p�BG�G�᪽��?�j+t�U+�]S��ܘ:�MR���Z�3���dd�P6^T�b�[ܩ��C��u�>��8���.��$>���|�m��*��S|�ߥ)�r8")�B↼8s�������V��9H�*"&!L�k/���A|�����^�Ȋ����È���7WE�U�]��/`�~zg)t���y��l���	]��g+șx0l+Jpu#��a�Y����Gg ue��҇;�S7b܁����HG��!�M7��<�S@ke2Տ�-O���p�3$���MJ��B����-[� �?aǪb~j�w1�ĠV�N���Ë�>����OU6�ޓ*��::���5Sú�a˲9�Ȱ��^������,�î�KŃ�=*�����8	��^�N/�CV�$0��$�-�u���3��L�T��*�~���x9P�{ﱅ��)�:����!��|��9.-�I�0SUŶU�&J֜t�-ݙ�ӥ���v	^DKG�a�r��<S� W����7�I����Zv��D�E��/s�Y5K��-�~+�����Nc
��?�q��A`2��)n+Y%�*l��Ahݑ$GJ� i=���4���	��f�2�j1��9WJzBcN���ѹ�W!ʌ���ts��ʨ��5�J�D��!4��T���޸�9|��+��Nn�fz�<b��?A(��j|-Yf�_Au�i�ܾ�;;<_"rz"�=�t�t������{���z��W��Nh}�;����B�]Wu�8u���,ފf]�l�S�HH�A59�z
s.9�h?ͶK���.|~��*դ�3�^�Fdt�_J{�J&-��\mI�P���������_�n2���/��~y�*�`�*�dU��y��tEAf �`ͰE3?VW���b�VD���� a�M~�R2J�Tp���֫���GM�v�G���?q}��m,���/7�EQs�\���,��*��3��H�Xk�S�� �-a}^�&�HI� �ҵk&�r�;W����\E�*~������C��@T���u����SM�#�^x�� �Z�@T(�_�\=.�Fd5%�ў���4����0�; 3fX'S�b0?�|��` .$��|:�}�X'Ń6�����iD�|�<�0��f�;c/�|Va����v����ɏ��C��f��a��w-��8!�i��6��B6������}Q(PbŠC"�ͩ%%F�2��m�C('��C7'U�2�Lˇz=�j�@�sC��WC��P��g�iU�7�kw�(啙�C�?�Ñ�E�7R 0[�����ٯ�b�]������R[�(})S��Cj�'�l��&.|0�99�R3<��W���_�jǯ�.��Ӈ8��I�p!2uEpʧ?�Ɓ�#C��.,��|�,�W Z+�?T�ڈɆQsG�34Z�Q��)�Rl��3\S�r��ӂ�isG��Ig�T+��_�[*�ke8��-���q$�m�nw
����% ��BQ�0��]|�n��i���qe0���im��}���p7j�"QY�a;ěG D��]`'��c;��[�3�'XM	��9�=W9Q@A��5'�JEMz'n(�\t��3I�M��҅cHЕ�f���7�5��1�'X���������<�U�-k��3ݶ+�S�O��>U	��%��T/����j�o�����r"rK~�飞��P�f������<�fƜvµ��n���z�s,��J�Q]q���}�G}���%����9 ~����A[#�{�9d�'��?52}����T�}ww%M��Ӄ�U5NEHµ���Ě��x���d��W�`�"�>hSv��F������VU0t`�'��rHQ�b���R���t�3.�i�͞^�����Z���s~z��
|ɱ���G杕&�5��Ie��%��/��gb��C8�izI>��F��k�B'Y ��{y�sC)��j�]��z"��ϲ���겷b	�W�z;?HƟ֛�7n���x^��D(,'`e^�SL+���}�u�U�	�_fx0�x��з�o�����sG�!���]r�h{��v<���ǋ����
��%,[�`a�8'�H�ȍ�i�1��ͺ�[eUS���e��3a"Ȧ&lso���7�� 4��mS^�)���K�(�R�"aمP��iy��{b�+��|�{���� ��Y�3K:��O�ČŽ�����-�Z\�,p��\�i���W��[`.,��dR6�՗KjrM|�XZ�Cug�I��o�Xy'�]��C����G:֌��M$�҃Mɗރ"����_j\	�.,ctE����%�B�4HP[��G���k�;%�7��Z���� xv%�5�};DH���a8DQ�ub�	�������`�%A>��Z��旾�V�	��,�l���Q��A�k��%1�E+����Z�4�����Ǖ�p�hf������Iz���1�����Y�{���-de��ھ|m�����n22�Ï1�ݒ�������R9���;,�h3I�8��Ae?�NI�0�,��V6�m�hR0�y��H�����?r�hXD��گ	��>B�3��*L�ha5[�vzp����4����y���DQy ���cpMU|Ilhl�U1Qm�Ⱦi���t&IaE*� �<W�?�3���%��'���{�e>W�/���[��w��Oq�l�t��^f�ʛX����/�n����=���Y�A�&e��VRO�3#E�r�n1�s�bD�u�����S�e�j� 7�n[Xۊ���������M+�v�>�=BHC\�]K���ni�Eb��ZB�٩n�ϥ#�瓻-1���aZ����Jʴo�>)bOŦ9G���P=]����R�K�IѤ�-ViS8�[��=`�0&Dpb���]HT
��g%�EbV�gt4��B�1J���<s;o��S���G`����O�s��x*�/��5I�\C���8��1(�X&R�1�?�O>_wQ� y��e���;�T/�U�F�24��/��ۼhWm�&Z��K(z���C�o�A��ߓ�J@j�|^��i�I-�-嫯��{�e�JS�h�hOT4d\�/����퍟��W��a�x� �� �A�3�������dX�.-���!E9���՛�ƽ�VFo�ջ�px�d�y�(#}���F�1��5j�}�d���%vl��ɹ�CW�
�{hZJS�V�2�i�	�o��/Wg�j�(9ʰ�+���	���O�*#n��O��[��Fx�yӮ��MX��Y�(��ۃ���hgn^��!�%D#s�p���ы�� B�o�tէ��������,��
�j�=�W�Tp]B��ĝ��b�$+��1���1�,����)ݾ�ؿR�T�`j$���h���~��<	���/�Ř�b `�Z��s�n�~w��1Af�?d�*���yf4p�!�j=h`h�4��	���X�`�E*��hKڭ�*�f#�0+¡g��n�Yc���-�?���F�M F+��y���_!;Wzy��S.��L�o��Q}g��DI���MQ�X �wS\���xd��ĕP?��P*�-"�X)��"j���v|�ʼs`|��n��D^�L�hr�N6�H����V�������Z��vxŎU���x��'��˧�06�f�.�`�"��L����
}�*�;$ �ꖖ�j C;T_�RK����ErZ�4�w(�n��D�����?�t1�$x<�K�K�.iJ�~�7A�΂��K�`.|d8��u9��Иmk��i�PD�����PU*J��aJ����=�F��tF���Z��O8������9�݆˻��[� �B�h�<�na����{���J
7��\d�R�3�x����ؼ�����!&���>N̓��������jG�(�uZr���$�q��'�7E���A���1��w���GѤXf������.4������U���(h��dGh5ÚR�?����ϱ��Jf��cd"�@fk�c�	r����I�h:�3
}�]�qiڮ1h��O#N������2	�p?Wޕ�#�	��g��I|J�ƀA�Cmj67�X��?O�Q'��5�S���yK��O\2e��|�
:NUN�Tǹ�D���x������T�>�0WQg���=?.��2�K8 ��b����+ى��\z���]B��&�e��M�����|�rVX���~u0j�8��ۤ���W��*F�i�*�YUEpS�#%��3�ї[���HI�8B:&O�g�V���z�C�T#a�g{Ż�k��Q1�P�(}5�4��{b?:?��-�(�!�ފ�&}�ݯ�e��ݕ���/���_��>���7_h��A%+�j{�#psTC�S���Y-q����tY��ԞJ�������H������^��S��ٻ����k�΍�Tk�����6-c��ͮ�����d\�S��(Op;��a�dnB�:��E�-�3[iң��v-`֘P�)�� T��	��`rZY�4�~*mW,+�0�� �n�PՎT* ��<q�Y�+a}�eƷ���k��2�˶�%f�:�ڎ�Pi��?f��2��>f�����o�#���ɠ�9d�㕉L1Rc�r
[.��K�=���v{�#.w���� �/l�ze��s)���]U7�\Km�H�"�v0uZ�M6� c$�AX��Y�p��=	���x��}���gy,9�������ε�T�x*���1z��(�׽!a)�7��h�T�����D��X��A�
��O&F<�@�~�Ϧ\,-8��W� ��2+#��rC�W@#�ϊ��:��Y�=k^��.��*1�8�tn�4i�T�.�!��R�F���)����D���sb��:����C����&�@sO����;(qj����yT=�����Rl�[��^��.�rZ"H�ە�92��U>�u���M��Wx���k�zG����B�g6�ڈ�r�]ϔ&8W�&��o�<�8�=h��C#+"��s7��bB�/�6ɏ��r�S��C�־}���]���5�k�ؿ10~�2:���J.]t����u,��fKz?�W�e��x%]�����r�|�'%���N�?B��2KC���0�J�7���FB���ak u;#���)���� X��LT�+]��%�k8�V������[yēbBs��C��[�t@t�]p��G�$+s��M����;uD5�tl\�}�W����\���K����G������>^� 8��"�ϤǦ`��QH7��C�ttc&5�7���$�#��X���.u~땗�H$��� �H*��6��TC�9Ҕp?3@�V�;<�^ ��\W��+Q�g,4gC�D�����u̠&�a��!#e�щ.)b���%�Hk7�Y!{ӣ�qd��w�샓�������g�Z�3C�g�C�q�(O������ez*)����Rr3&W�p� -?�E��'��t���u��7�lI!BsB�.G�V dzP�ySDMkh*VEyG�z��K_gtbMPJ���h~���?/u�P�K� ��gM(���7�&�=q�W��ٖB��+S�°�-��7J�>����.<'�M�����rD 䫫d��H���=6�]����d"}���T��d.�s�����G9�~�1u��Tne�ВNy:;$H�Jlr�hЊ��<��W�!-�d��>�=�S�9+Y�pd��]�}0�햃SU�B&D���:lk6@�7n?�w���{���+��J�Tx�D���|�t!�Z�p_C�@�qP^[A�oB�oJ�qUk���T�9��,`�M���܊���ڤR�̱���E���1y�1�K�u�M>�myK���Tk8�Lu������4���n(��l��ew]�g�2���4l�OmHd���A�ڒB#�����V�ـc3�c\Y� ���#}Z��Jbr���+�m�U��4�=j���u���hG������*|�=��/j�-տ1AHH�����C=[���T}�j�t��Cy?�3�ڝ���rs2=X�k���GuMˈ�ou�N�gބϞ0i	��v����^7u[�g�Z0B�gʩ���rM��^�:��������ܛXc���ݤA����M%h�>\����CoYb+΀XK)��ׅ2I@���o���O}�"V=�Y��t���7 �����do�fΤ&?o�����S��u�<�����2�;���>�	k�C��}G�S�\�>+��I���+���O`���x���%1�g!����`�J�r����$]ɤ�â�?/�yr(#ȕs:�-���8c�r�>�V�{^C�9�7B�HJ��&�0��__��4p<*/m�5�������p��\)��6�#�����T����/�)�d���k�%��׹@�	�q��B����G�k���d���~T�T�MI���E{�
�*�� �e����t=f�.z�'��=��m����m`c仭>ʼ����C�Z�\v�x	��{�"	�J:f�Kk�Ю��ɻ2�1E��;:��)|Z�2W)�M[��-I�$��[Y�J�IN��i�+�d�������<7�M���ǔ����@����?:j�+k�?R�MƲ�C�;�s#\��ժs�);�gK}�tC�f��g� �ɐ���p�`��䀅���W>���	C���X���� 4�x���˃UH�`�F������ىs��BT��д	�Z��8������$��X6ְQM�X���/�4��	X���)C�/?��f��憃�Z����E��I�f�N�2p�rn�Kz����+J�۱�S�]ɐ����c>�v�鬵����X&(M��%�^gR����2�8�fY����nf���=�b��!ο�p �p�Q�& ���(&9�:b�1>�R�Mn:bVk���U���)��q�`� ��D/�a��ĉ�$��x:�I[$��?���o2ɞ>��;\�l���Xy�u����C8��� c�IϜ��x�:8��l�2��]L�h��i��1#�"�������T6Rf�d 2Ȩ��Ty�����4v��m��|�z���c2r��N���-�?6l�>�h��� |o�v��t�z%B 庴�ut���g�RjA\f�w�f?\���Msɾ������?�N��Y����%�Q��b��lD�$�*�^r��%̃zg
].��-Ó^��`��W�ٺ5H#ŞW��E�D�쓓?�F"�x���K�1�^�[0[��Yw���0s^J>ȿ:&���7�G���jϘ�I�#c�ibu`;n_ky��M�`�;7���#�o����!Gg&��AM������՚_�8m� E��~��?a"�4�l�	�~��/l8��l8�Wc?�H�H#�r��轛}L=�^�/���ܵ�lD�k�]������\
�UIX�ؿD��S۰/�O��n�}����oQ�j�9v�D�c/C���_Q/ MlC���!T�s��t�' j��<b���QD���ȁ���Q�N!�	O�1C��	�f$���1��,Ӈ!��6�}M�>�0��ʌ�	2��]�5	ǉ�-W�F�I�Ɂ|Ag�3e`�}S��S�0�S �u��к��|�������mr�94?%_��\�"c��OG2�����6z�[ u8��2��8�$��8�D����=�P��X'�̱��am��}���f����P(�N��ت,2g8j`��V����Ш�(%G���J���ְJ�O`7�O|�+Ofa9�^clX�,�3D�X߉��v(l���Z�A'�0�D��y�5����M������ڴ�D�լ������\�՗vmjw�2eޣE'��taP?%:`�0�5Bľ�J}V�E�}�}-_о��K�X�,�����؍(��.	󩞿bۨ���2ү��1Y�1O9�Mĵe��-˟��Z��7�����w#,%��('n&���i���`5�����K��L)�'4w�V�#
�hz���|�ޱ�TH#0a)A�mY�2�'�3�**���a��9b�0'*~�j��PKMN-�T�.��q��:��Y�@�q��i�]=����f�ۭCK�����^�rwz>�M���9�3�Գ�`��3яD�j����S��9U7O=ǹu�H�ŏ-� ����?���:8���pE�����v_��@��/JO48)�sX��8g��ې�_�ק���dS���|�)�Y1]a����Z)��T9���%���|2|���P���4�5�>��0�n܈Ԍ?5I)|�A�-4�[l6Qc�F~eϊv�E���m�=cW/�������;[�2�<P������v���rػ�/��~Q�A5��@�Wp?��hc���� m�\u�0��K5�7V	�MC�N��v˕�N�.�6�>"����o�&�βo}�]v�eu�+:��
N��lئ��)1��Im���j��!Gਘ�_i݇^<�V�"�h�@"������٥$9�T�&^鸰��S�iv� 
�L�ө���|�BF�T?f���k?[�?��к������;9h��]R��\U!��ɋ)�e�� T��l&Fw7��!Ȝ���nWtA�n����S<E3ʱFi(N6(�u5co��T7���_�g}�W��^3 ��,�>V������_e!j���ؑ�*� !CliпFyo@ꤰ��C��8{&��׿z�r������T��g�8������>�6�$.��ř� �V�R�{�#ԗSl���D�e���q�v�ζ�6��Y���0H���ȫGEa$<s3Nol�SR2�v�@q�oI$��cU������Bc���-���+!\m���;y3C֋��P���Kז\�jj�1z��LU��E��oR[���3��H�;�}�jj�W�C��Kx|Mu�n����ׅ@��J�p��}K���M�!)}΍ewë)�CY<b����(p���&���)h,�]��I&���c^�)��l�`>�;�ܶ��L}��̟?G�$�߂��ώ��/��������詽���l^��&�S+n�Q�u�7(m�x�,�_��y7KDC ���6s-���Mޒ���N�l��M�l.�����.����%�%��k-u� *т�V�5q�J�k��+O���w,R캑��zU�o�f3�����������yV���tf���qQf��.d lOH�b���o
�j�b�o8γW�a��gX�Z�^�����
9�G�G~}�b�	��ռ��Z-@HB D`����S;�%cшk^x��K����J�e�%OS�
<�V'<��K�(�a+�����:����
� ��y�rw$��>.�Ϫ�;3^(�0����� �6��3����8�/-ľ������n�m�>v�ejc������`�u'��ͳ�Y��G�Vy�S���P���^��-�,�J5�Dd�	�5��^�x��7���!�����n�n�C
i釒{��]�����D�u�0����-؞l��p?vbwJd�(¹,`o+����c�w�0�D�<W�(�F.Җqm�UDʿB}S� JFL(}����q�{e[�>�`@~Y�$x 2K�J���c�z�H�"OTᵰ�AɍZ=s1������q1n�IrN��mJ
��ǒ�҈��P�:������_�X��1������3���h�YSe��� Ֆ�}&TR; ���~o�37�k����/����Ξ�]\H���J� 6g@�.������] �Bv�5����y���E�Ì��ץ�������~���cm1A�� R�[O�HPMF�$KP(��3���"9[b�������cW,�0�Kw0�ś&,��|dl�����1$��`n ��2�Ч�
գ	�m|#"��`�' ���s	��9�;�[a��wI[�yL#������x�M��^���Ug#�
�qBe�^�\e������ꖟy P�׮�!c��Y<�v�?�g|�o턏�i�^3^��[���D�#tn�'���s+h��>��7�z�s�G,����R Ol��7�x�K�U��<��&Jt��qNԸ����%B��(����`Z��f���lS
���'��a�o�s�{>l'�HG�zV�����5�-���n�+{[�߲~s7���|�hN�U��>  H֗B�JUኑ����m6�Xlg�뤏��,�S2J�b�@�j��!�Rb��4����z$2��d�����I���y_�������ik���!͂?� �`�Ha�90z�N�&ʱK�{B��Y��Tj��Zs�Kz��I;%l\�����~��
Q����U�ik2�;oB��U9;p�2�w�I�o-V�Ũ^��&�<�લ������-[bZE������e�rG��?/,XіJ1WV�ƀ��p1��':%r��@��'w
GW���5���m���� r�T&1j���������"���� 6WRT���C�Zw&x{��&��m��5����T1Q/+9�x�[�(��6�b�����y��w�,T��R0H��Ʈ�Ɲ4dt�~]�*�Ly��)0HC\1��w�.���.�}5�!݌�q�;�;�cA]���8�k�#����~��@s�!�M�������^Q�> p�!�A�h×G�oW��/�qyн6,����~Dk6���U��x�0<����_X0�ڦeK���[{%{+�Wr!�~z79ִ3�f���.P��9���
R��`��6�m'�3}ٜ&�[���п	�Z͆\�'��}?�q�4=͹ee" h
Qb��Y1���-11�' jdJ8�9,d.X5�Mk8 �-����I��΢�4D5�c�5]�o�7wqg	3zD����(�i��I�9�F�Ɗ&ηŵj��Uk��x��30�f��i3?���,(W�0���u����麄N� ��(��-�H{-"�LX��[�$M�"u[�ǋ8��Q?A7�P��P�a���z!bOu�g����L��4���V��s��F�'S
q'�1�N�I[(i��4-O"��jWwE�Ry�̾��qy�{]{W�uH9��=.���8���x{n�nMQ�B���5*[��7!�dR�{n�!��+_�A`tg�C�2uצ˃���-��|im��7qC`�R�b��q�ox�u�aͣ��_��|����/��/�c����,�v&�s�lU��r��g
Vt��,N���}#\��G���������=9�S��3����e ���@��1�w��r�_{҅9���U���Wl�V�*�l_�ίį�yɅo9�(���W��D0vI�>�k�|~�V� ��k�J����Y;Qn��D�3�7�]�;OTy��wP��"?R���O��(�� ���1��8.�>3����B��28�":��ZXCIĝ�� ����\O3|uq����/��*z�}�%��8��uo#���<P�|Xm�n)����䑥����0:˼�������w!쵲��W8�{(!��\���&����Ex������w��i2�,6�bV#!\�j5�5V�q��M���Y#^�{�d^4�e��bښ�������k�0�c� /�0��t��o�K�ti!n�r#���)+��v�ƹ�aW����\Y�hC!����І��AO}���kU�*�)'ҩ�[����������9�ڡ�]>�mxQ/㎉Ԣ[!�t��i�C�-�܇.t�(t:j�k�	.�f�P�V�g��;�7�t������'��»�׍�����6�2x]&�0x���c�O��o�
{5��	Bu��V���,����鏅�b�|�z�%���fߘ�Jfs��X��N���#�ߢr/񩾤N���^��h`!w�+:��i.�E�4�q��q`�b���9]od,��M�����k(�����N�z�R.3�Ipy��qU������& !Uv�F�p�X&��+`s)��l��T�t�Ƕ�������*��J=���8��H�-��c:\q:�bA1$����0�bm�h֏���/b��k���f[=�?*��߾k��9 �&5��|��

Mi��L@�����PW�Λ����g�r�'� �����2�c(ҫ#��8�)�#,�\̖lrx<I�Xs�7��G��B�)=��#~���F�an��oH���X�����p�w#"v��	՞�Y��~�{ |�T�����$Ư����:����@��-�ի �ԓ��E��Ub���'G�'��s�;n��[�6=���џ���c�Ջ�K~��}䪽���ǚ�STx�E'D�k�C\��h����܀�9KsN��}�š��v�V"sҡ�������� F�S�ɔf_E,NK�6��;�e4��e�/�,a}4�aHӗ�O>=l�#@����%p�=�K���n4����0�&���Va�o��.�����N�U�L�	���J��X��q�P��?�ϒ�E����a�A�m�us?�r�r;� �HMR޼��jMV����DD�֚��	v�oUz@�^��'L˔ߌ��<��9�UUb6������zΌ��<�%`]�꾇T����2�fR[�\!D�����؄�xv�;Q�Nd� �!W/�WKǣ�u�M+�XD�W���>�Qˎ.��g�Ņ��m�J7
)>-Mv}.L�i'�mO-��TL��n��yD��]K��k���ˈ"���8y�u���U�ʹ�3}�iK��g)S0K<&b�/�Z���M�xYI�p��j?z���d|�wp���\��=;x}��A>�#;M�Ά�)�pCb�JA������[�(w2j*t8� ��@$�~r	�����ϴ5����@d���;ϯ t��!;�8M%k���9 @�Z���^n����)sYg�jQ7�/6dx�a��i6ݬV�­�aG怏��[�߈FE$�/k�5*�| �~'���Z��È�d��2F�4z����Rgo�㎵8p?�T�н���+��`B�a	fC�}�딄b�`S*������ E�n�VV�W����+\�+�,"��Cq ��5Zz
��Y�q ]�����f�6D�Hnp��9e>���4//�&�/&��� &��x�1��{����b�`Dy��l���o��0�9�w21
�z�L�c�-
e��W��yѭD�U5Q�ި�K���]v��K�
�A�x�+�ot�g[�f����4�$�lW?���jv��A>2sxj�VZk���!��Ȇ����;j��-Ґ�ǔ�4IG������V
�}Oη�!1/������3�˔ ���z4^k����..���k���*�3�kv�t�I�f�[��,eS8H�2m��U�"H��aS!"sU�+�al�Wg��"���<�(�<�V H�{,�/�7� Ka~m�j�$z`{V}��^O1���#����mk��[�+�y�ټqL�~[��%��x
@X&�p���\5�-��=_`�Y�6�ǅ��d�����b+U����Wn��qϮ7&��ߊd���{_������I��;`�b��R���"�04������N~�5�G\CU9�7��-��CiE�x�a|D�!�&�7���^�mb
�v��Ї��ك[Lڮz��X����_��,*"�!o&��U�B�b�-κu�tA��3J!e���/�F0N�_��pΘi���E��я��6��[V����X'n�6�=���a� Z�]LCCg�?sPj�!��3)�yY�4����"�f��u$x�,���?��4ǐb#~4?	���n�?�c��,�2��IIݦ�:f�)�B�?@Њ�9����[�Bxh���5���"���O��j�>���5e�s�.W5��AGuJ(**���n�~��2�_x�q=��#�����z�l�75��9����p���3v�����O #�Y��u~U����Џ�� �	my�QrMM��)��M�G�+r#�̝�Q��)���F�~�yT��O��5�Ia��� ��.@�`£�os�D�wI��5'����Z.���u��F���fW�9�fT�6.1g�bV����P�P���
(���r�!!�`�Uɹ�*p�����4"����țk�r���Z��<��`�a�*���KD����M]b�5�g�/������Ĕ�sP�����'��3�υ?]��[��V4�B�#���
�/y�H��\�RE�?!��n����x��_%!Ҫ�Ƕ�D�l�=�#y3'�����"Yo17U����Pa�[,��g�gP�ev
�E�{`�O��0B�hb��(�r*\Y��i��l�K�}OE�qw���|�;�R�����; (w�p�s{�r��e4\*I�`Ȯ���'e�U�E��w�Kс)Q���	��R��пݽʁ��	0���R-�a�4��<��>��b+����l����"|�0����c�IϞq��ܘ }����ߐ2X�rh���ц�Z������Y���̄hD����W���=n+�PԊ��8�`�ɑ��GA��)���EAO*姛��~�O�4Cc].6��O��L�Zi9c������M"8��s�8�}�t	~�3�.-v��iS���JS�?���r�V�H�Q��XnoB';�?��&	H=��k�*$�Y���t�*�0j��k�
>����i���k;V�3�}���D�vc����Lze��#����E-��vk���1dy�s`3] �-�L�0��d#�������0Q��`�S,��8��������s��ď��j�x\<r+��qh���p6����T@32j ������|��J��)���
�͓��Ϗ���#�߉��L?_^������U��!W�q"B����яx6/�*C�eT >�� �D���Kؤ;��J����T��b����D�58�KQ��.��Lv	-�6U��4:GK��1�UJF��ӽv�H�'�~Dp^eR96j?��<���Mm��O7Q�eS�wn�Ӳ]���KG��;�N���B=�2�#:��^�8��E�z �l��>Y�O�ś�̀7~K��^x�8�F$�v�^׵�RAʙ��@��HB�ub�ʣ�D��C�t���O~R�Ǌ}���U��N�6�Qi3c��D�6�b��]>�r8���SkS�}��!���_��`���b
�|g�ӥS��f��s-��6�:T^4��H!��TN�ܲ�a�����X�� .e
���(�������F�C����!hb�WY�������[�C͠�&FM�^MI��`?Y{=�&p/""CXpum�U:#��I��ŐKR��=tqʕqj͌��u��9��J����)""��P2��.hH�g��
�@�$�$wK�{��sS��D����tViV��dl����aBv.��T��U�;h��R�V����t8p� �bW	�f��3�x���"��~C6vb��j�%1����Hb��v�Vػ6�^G�RH_���N�m����G��S�����������j�+
�n�<��d��)�M�Z@��9V��"����P���om����w��z��&���l��6���'����HrLu�&x��u����; �� ���S�y3��8�#�y+g2J
\�V)����\N�3~;m\�����
D:���&�/s)ެ?~��"�ʻ_��t�_\Z�������s���r�� ;'5��!yB�r���(�ZiJ�56k��������<XJ���勚�Ǟ�`-ּ���awX)��-�?r_��\�p�KTk�D��ݿD���c���1�!��a@'��{U�K��5�GȨPA��2�G��5EɈ�7�p�G(`T�S��T�6��w������s�~��T��֨��݇����얛� ����Q%�*#�9�OFc�f%���I}xb��4U_o�)m��c~Jr�7�g}�%Gwh��Z'��q��&p���,�P�Tq��2�b�G�n�ݱg�kΓ{�	@�zT���yj����`u��y$���_�"Z�m]P(UkQ�u9l��g�!�n�`?
0�D�j��p�%7�]� ]2�x�&$O~<��>cV)�iaSW�E�RH9�䃻�2�6�o�H�"�p�_�X�$�sŦ�W$�$ʶb�����΁�6�x�AmIq6~_mP1<��Nh��tZ�We�Kr���MɼC��#�_p��w�N�儩>l��~�8���S|1MrcHv�2��'�9�?Rf��%$�_�z�2˾lv�����O�����l��KEF? C_Ԝ��"܄(��)�}pz��I�R;�E<��jO�W�4��gvRH��,�C9�������:K4�Q)�|�������7z �;m4��7MC�@����A��t�wHO$�a��h0����1]������k�ʝ @o\1��� ��tٷe��eV�$��$;���W��^N?�����5S	�A�:m�Ց��qK�V�^>��*�h���?�� &z K���L�)#����-�2�oC�FG\"4j7�Do�=�8���}��i0���d!�c����z�>��j�Aڻ�;�g�)<t��F����0e�S�Q�י%�x�����4<Je���r�fN�Z/l0�2[XJ����=�[��:a?�YS�Ք.+XdMc}�t�|m�b�U��P�9�=����ԞJ��ղ��@f��s�@�4���B�������^Y�=�%�q�hq�+�i�������@v�_�^��D"��}� �w����D�[�������J��A8ʵ4̌����'1~>z�*�঴����T��;�d�_j��Z�9Ȩ���a�%_z���fwP��֦2�˺� ��9��Z���0@x0��䈢�G�Y����s'���f��{_�@"�:�r�WZ���*������^h���˩��+k�.����1f�XB�i�t*��t�b�>��&T������jה��{.�K����P�.��	�s�p���-�k��I%�+�/R���/[�O�¨������X��������JMR�$�����v�u%�j�m�x�Ԕ"!��,��@�P��+�@��E�D�\}��b�C����"	bE���Ӓ���x?�N����}���t�m:�1<��C�v���[�$d���t�0U��'%: !�ѯ5�P4Qe��R�����a�ˉ.�km��`H�4���dHhxp����ql/���@�����x�w�:(��0	��G���7ũg	�6R�2v]C��{Q>~Ĭsp��$�P�D�q�P�`W�F�J�s5b
�, |�bL�J3:q!<3կ���9I��K2���D��q��>�\���i#�[\�RK��}Nǐ�	�"Cz�4g�6��ZYǚ�M��^���%�����Z�А	ZU}g��w6��N��ҹ�T���iQsnC���吝֢;y�-E�{���̺.��k'gM(���l�/�������Hl�>�����4]�4qN"��sW���������X��D٠y��g
��E��d�Z��o��n�O�J:�y`Xx6�Od.�i	��}��]��?�՞����u����`�qf�SY٣��<����=�]G��u��k (N�LK$e���m����ջ�ڴ��.u#�>��L��'?{�c�#O6&ȼ�����)qu�Hc�{��C�&7�z��̨�
c�kI��T�T">׿k���P�d}���>cZ���D_��j����!g.��騈э�,�� �Ss���SG|��M�D3J����	f�����l�	�F�ڧ%�4�y"<���s�8.�hUp��`S�uYE���1G��f&w*�䴻�uk
�5y�c��� Q�Bw�1l&s.��jM�26�:Z�������,=���	W̏��g��p��l��e`�[h�Im��-�e^!�W�(~�c�{��m���j������!��Mk^�ZPn퇱�2	T�y��4LD��x��<�%Α�M���G���(� ��^���d���p[c/,��h�	�eQޥ1�2k �T�:�E���l�'OL�U[r��F���-�����@xV���38�>�����B���-t�ֶ�m�3�a<�Ā����t�kĚ��Ō �1�)�N�צ���z�/���4OF�k\�G	�g`]�f:�}�%Ԡ)��w���>�}�����z	�����P}L�oYŌ)[Aс����EMac�|f��dv��z(�SXJ9�V��?M�V%� �Ҏ�ٌ�&a$��$n�m����[qR@�8l�H"B3Ep2�7x�Q,&����4�E����cM�P-b��8�t���j}A��0Ș`f�3S�+���g)�wg�p�gߒT��{Q��7�b��{����,"L�(�?��V���_�B�ڦ:6>�W;�+0�t������`�Ή��mG��Y�X:��ִl���`mq���-F��70�ς����Xר���"��	�9���a��Q�+���ukQ^�Gnk�����̝exM��k�Iک������CNb ݋���[���0\{X��7?W������dW�w�8L���=�;m�|H:XP��v{%����U� �Y H���}��P��:hEŢ$kC���5>��'��c�$�}��&qR���0�u!6�O�T~��5�XY��E�t̐`�0}Թ,��'�(ʿ'й����5.5��DK����� x?�=<W������~rg0� sX�����j���Iz;p�
O�{+��s�]��;sE��L��עA���6(P{�,s��[�;:\Ew��j�~�>�?e�'"b����gS���b���[ٿ���i �1�,9l�N���z	~a+�bA&�@j9E��]q����Y�j{ņMk�����ȋ�/	h�W.[?�Z~#�Ab�B����?��Z����ʐ�װ�qeu:�~��v���
ALX���i���	���6;�V��&�E�X��R�ڣ�a+�U�%�ٽ7OMo������N!ƌ��(7`�H�'���l�T�Ӗ�����T~�q��7�{.���3�9j���H��p���ܝ��ͭ�����$�m��v�*�Yf�J��#���q�T��J��=z��F��e����"�|uQ��hMdG��:����/"tk�������O���O��f��,�8C�m�]=��'�i����; G�WKD��2G(�>J�K��c;�(Q��U�[����֏�[�c\L���]l	O�px���;����X�t�����m�6��Wۯ@&��/n/��vmhc��TG� �������F�'
C{9�������۴���3��]Yލp'�m��X��Z�O!�:8�P�s��o�Iʳ�.a�����U'������lr,�[$�`*!�5��X-����H�=���J*J�Q�z�p�9�O/�ݮ��`��Kk��!����ң��SceU���Bh��^��f�t�E�Dk��05ݿ�˱� ���ޱ��Rh���Ѐ�y@Ђ���v��6�F��bR/�*������DW��CiS���y�w� 5k�#8�6�#u I��r�(?dl:/�.�tn�;�0�wa����@���RXA�1'�	��MM���*�t�M�� �5`򼪁���&�5���ȪѸ�0�������"!ζn�z�)	e����� t`ܯ�DǯWA���!|.?���cvTi��T@wfd�y����/~��|YPF�e!K��Ϯ#$![���_jD\���b�b�`覨
���Z����&܂xZ����R�-�ȟ��|���hU����ܪ���xg������,��WC8#��<�V�`���|&o"U*�Y^�}<��pQ��%��n�; ]��4)�C'X#����8�M!��&S��F+;P��e��Kw,2l��"P]� ��K�DAy������}Oy%��Q��,��G����ě ��8�Z��#��~�|�$,�VUF��%D4��S��-hp��,�\.a���L����T�=�j�;E�\ٔ,g2��\v��'~�)§�e
z=�X�/���~z*ҮW0��<X@���تT]8�'�C=�D*�?����s��$���t�ro�ZVm�����pD����@��.��ʏVT[���+��������K�ޱ�fVk���aO�C �;��_�BX��7&���}Op�o���N���}<��PM���{�5��zJ�/�)1�:���]!��.��b/>�j�ȧ�5�>�wj��(�9�2&�96�|Yr�qi�ۧCW�#���b�Ep�o`i#�l�[�S�?�X�%
�<�����8?�(�x���W�O��j���9}�l��\S�}���V�-]�$�v��[�ߴʋ��V3�)5/���*�F5����oz^�H�GD��F�A��@��$��+xXn��U L�0��J�!!P��~_��_���P,�W��~�]�t�\����a��K� ,a�܄�`�������jكdKx�]�޲k,D�lUDw��SB�l�Pɨ"x��F�a�ͥR�ҀvtQm�d��Lwj���d_��D���"𰏌~��q��.������w��M�%1G �?>8�58s@��)��܎����(�)�K�O��yH��TF� I�Bj��=3��ۯ�|#�YD�_� O�~���xG�#Zt�=FYm�,H��p>���1��v�e��*�ZU\�nΉY�<y�:'ǋ���\!����'�!�> ���
 [<�
�:w��ޥ2|�g𽬏ȴ�`�XŀH7	�F����) 6�X�J��ηk�UCL�R�ګ�VIrֶ�3	�������ظ��=�Go��������j�Y�ǂѥ�-��d�D�mF]��"�A�o��Aܗt��f?��r��n��}��}�^TK��@� e�5�]�h\�Rڄ>z�ʇ�V�G���h�� ͐���YXNa���܉a�4AO�U����Oc5`�RPѧ�B��Fe��x����\X�f?Ȣ~=�AR��H��C$8hM+��Yz~����A��P9���+���	�J)��UD-W*n���uK.3W:�OrО��%�{�$�5�v"��7}���ɩ@���h�^�!>��g�
��i�yo��c1�f��Z{�L8e��h�k(�C+���ry8u�#j���@��m�-����Ȏqy%��#~NK=�U~1(�_/�TRk�́l5�B"?-��CR1��9�5���9�������Z���X�#4�MV+�8ԯ�xa�ót=7�O1l�}�Qr��ѩ��*�,6;ܝe�	��jj,�> b��d~�6XE�;�`]�I�d�� �����-lC�ʦ8.Zp�ʊ���6�V9�9�N��3l)d=z���+س�{"�~�9�����M��<��@�(a���Cܾe��FW@֣SΙ::�̋��i��=�HM���NS��Z�@���t�c�p�*յ�Q�܅�i!�5�qt��K<.��R�u�[��3t�g��Cz�����6G��EF��$3�Znn/��{Z�FZc'�Ю��R�����$�+�Q�4������r���vBv�=���*��ϖ�S0�C����v`�lMC p�6�6z.��KϡΙ�j�m��>���a?�\�������@%wq[�#o�s��e��2�l�D�닗��9���R0�@p��=�v�6Q����-c%+_
"�����z�	���r��u�q>�A��*S�٢�W�uy���vR@�S�*d��6�=x����m�T�ԥ d�	E(����C�c�H8U�J����_�~;h���? ��wW�Q�)���O]ߏK�(��}1�G�+=v��ں�����8tz-���q&�!Z<ˈ�<R�:�j5v�)Y��c����^DCUejFH��T���0������/���Y�?���X�g2�ɇ��m`�d���~�%P��)�@H驈���ur����$6E�T8@I��駝i�=7�Ӣ'&@J���ΕF�ˀ�:|K �*g��[߮�p�ވ��&1o ��_��f"~M*V�њC�"N��e�'��>�um� S�a�}!���n����b{}�\��L,��g��{�J?���0���Fdn1��8�DD<��
(g��>� �y@�P����y��3;>Ҽu��Fbh<_ؼN�gꇽ�:-���L����XKL����>�ܴ� ��D��"<5��E�ϟ&7iI�y`����oKҰ���m�!�����[�B�d�{�e���P� n��L�O�/�����U�������V��q?ʪz+,������T��`B^�d9;�[�Lk�b������;�%���N2b�n!z�7�y\c��c���V�JǠ�FGW탔"���
mz_	��V��0�O�
!��N%��*C�^5���xOtܻ�Ґ�z��'���G�=f��R�{0�Xu�6h��_�h�S>��F�K�䳖s#�( t���O4��W\�b�O�#���(�r�1��sܚ���gʃ8dv����f��V'V�J,�n�����e���6�|����q�COK@C��AG�x��x�2�v`A�;JI��+���E��\Fم��?�y8�@jLz�T���Rv�(��*�//�=���/e��Ʉd�n������K=��ox�BC:�r�t�s����|I����sT��/��N�k�5��"��"����gϚ�t�ǌw�R� �=Z�� ��4���C�l'��.aF�O��CΎ�/�|VbJ�q
҇0��b��A���}�;27��3��
"|�ez�uJFf�9�*�������s�n=c�El�?�R��}\u���F�)��_V*3����˽C�U�D�M� T$y����\fhs}�������-F:v���/�P]=_���	�m����7�ՈtD͌s�߬��ݨ�G��B�@[��+�Y�"}M��'�ɺ)��m����1���kgO�I;��1�4�"�X���e�\Y���cU��#���a�Fy�,�#Hq�P[h�l�hWEa[��tp��[��}(����Q<
��;z��լ�'?]0�+��)O�{s����cO�0c8[�g�1��_��>� ����7���4	�X�A��E��B8-��S�V���19XW�y /,8M6��z?�6��B$��W�9O��y����3a+��,���f%���/G�:+�ə�T����ƾ;;8�L:�(t�}@����Z)o���]>�3G�k��䅣a���ؔ��+,E�z�t�� B��cɜ&�鹻qY���VN	��Y��R����;'�����MH��]G`iP�*c�,����`��T4#�F�t6p��%W�x�tk����}�W&���U)Jw�:8�^ 
,�Sb��.介��FIQ���D�7p�gv
����~ܙ�/5�uv�8�ה�.O��]��ժ,x�~G�a%jV�f���0�_K}�i�}��-(F]Tz������E�	���z~/�{Kyz!9��B�� }φ�_6,b��r�КV<���0�G|������ξ�ʮ�ʬ���C��b��ƃ�I��{�f�,�z|y��:����	8��g�Z	s��&ZCi�^����&�5��Ks�thCi����NW�+�E�o.�&h�q�M�'6��M��5-<�H{%�A�J��%q����Ax�w�x��텞�lt��S����øS�0H�x<�c�p*��A��|z�v���/�T�ai�(K
I,�;{�3�^$0T�|�3��!B%ɽ�t�ߴ6m.7��?c-L�I�U�����ǟ�4��w�.�Hx�1��V����6z�U�_mS<��[��]	"��1��Q��K[k3�zDC��$�o��Ȩɜ�H+�bg�°���b|�
�o# �D�o��]_}]-Ew��Ni'gM���@���J�&����G��Z�J!g����{ݠ &�Gk�'"�>莝��.�H�9����(���3��6
*+c�wz��C�0��n�!_��w��$