// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Y75TNeOvcBU98TYhdqwntIAxdBAyGkYweAXYiyW2Z+4fVkBltEb9K+33/UT7GEBjRuDMh0zNgd3/
X7ibeobFwaxdSU+0GRBhs41C7q2BAi+KxnhjNV7gt/TjAdBLK04ItGI+spvSf09TjUHPrrI/P22d
8FabRkmWwgGjuPGIhrKAN4ScBOhQI1YwwJ5TqP5bvpKry2AftDT2lrTHguEKQBv14w0f6aNZwlbI
/FgGOW/C7H43hamKWJD32bvq6yAf59zs2ffmkSHw7fyRe1cHSevCBWIeXNcdOEUcoF88ySq7bVE0
lSvCNWA126vMvpATeqxenezerDjeq7j87/sXmw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12784)
jiBjmY5w650w9SiTh//dtyARWMAfecbqHPd1Vz7oslEGmHeQhc7TC2A3GGq+BO1JAHJdkLlOF073
c14cNSzTyXFOSte6QokFUwvrE1zd3qVR5BMFPD5Pck0ppXom22PILUyq0x+7TZIsLXgos6JOgxrj
EeEMEauakKOhLf9e1OFDTCXD7gNqKMBop+uzkC7ftOCQmpmZHYkv1WNnxEPs/nIJIi9RmqwHR6pE
5BckaR1ziwCJaBmjNXnnstemtdGNb66hRgVL8VvPM9GkhbgXVAH/K8kaby6WcTKIqbJnfm/CiQso
64LdC3eslj1Jdxrhzx4BcVHGsl2crQJ7go6AUdXoVl+osdVqN9weTye/W9y3QFaw+rda016l2PqQ
eJSPSXt1CpEQqRXEoMelr3l/MBVep3WxZ2bAiJj4CzC8FXKkFRGPPAsygaqW/0VKNa1rVOCv5elN
lPFbVWAUmjLGVgWAQbVCbT5QzL8V5x1r6dISh3YMPd4ZYkdR30+mPF/KLr8Agfkw9YPeOC2j7gFH
qr25GpFb+qk0QdY/aImgpVzfrjlF6BDp2CwY/8Ts3gmnZnkhGpZHP/b9/o97SbmkNc3KuJ3u3hAJ
UQe4bFlk5dmhqZLMiPN44LmRDGw3x7a5RMVXP+tpvkqeP/GViDgErrKbwUzrrfh9ZZFfrPb0s9LQ
udNdF2cl7/SiQf+BtqkceR2kj+hSHCcl84BOh19jUU5XmKwNhn85CmtBjygY5Zc08fJFXF/Cna9U
wc8YTVxPAY/cbs7OpX6++zMMP1mDBcQ43dHyNEIKOGSwPQ+vENfIwjyIteWcxqxgWtKetZSL3lC+
tfrhIdCZuIELSTnGD+VJA5xXwNZaz0glxJeWOYOX07XgaUl3qlHtWRQ7Lrl//N4NQb+aH4S383In
GhlB/q2cwPe6mPtHYtwhRkz1Lc5nELF3nuhgYNI0U1pbxmAOkWZp9iW6e0ukwUSYMGcFhnBg6xU2
KtEuB0cXXYVZMhnwT8BZSe65JmTSUta/931DBzbRsiEAC/0hoeNiIzhDknLaazWXBndJCz0QNUIU
qT5Uyoq0YK0tonfnGApAyS/BGix4xk7GYw94EeUz14JxLI7Mwr4I6ihON2/xV8zBCyGOKAaTGI5U
pg4OeJ4M6gNlqlptgj247DkKwHH4PcmM3X7Nzv4ZC6DLm+8I4M7LiRJgqlWLUExrhfInK8ISngbw
NL+JZMRbQRKoNSf2sfatoMk9VGs67nT7rSUIT3kcIwNcgJyUEBthOznQcZzqiZNYKD+ynaMKg67o
X4huELjYnMUGwoIOhOPZ7ndcsJV8+m4AYu/TueYEnfrQcFIfhJjOX7LSFtIRmK8cUqXi9rPRNWNi
M77XWfW00xDtJaG1lxDrPm7kOzwAPoMrOY3Fa3Q3sXT4fUUJi5dBWMlBM4klW7l/1E7Ih4SB+i4I
S6ERlstDolI2E4DKCmwPBBx9UWpRGGgY/0Wzq73WNhMBkwabMZms+ABAPOSj1GrDYbcYssfRuz9W
asorndQAwKMYSi7/sNSblh8jr+qtpC1H91ZYnvb81dYhab4E5v3tb7h+PqSEXLz7510udoV2Len2
9ZfgIarg6MC1EKV4Z+YKO3Y6w4Z+0MODGf/DbMxN9suchR+mRPEO0gaOEz3yaaNQ6iwNHcdsU6dC
ABkeN92QO1yqaKyWWRYP4pzAAAg2uQ6DUixXJwFCA1zc2tEGxO33jKuf/HeX9le7zHIluBE0j9kW
Jqz6j/onogBaUa2obIdMM5LxQ5MKO3KJJOPxDunyVv3N6SsbJttpXhQ/tz9vwMkGZE1tjoXowyji
kABsojsVTqymnMbF4J91tVT05Nc55xfq6+GoEzS4QmeMpJ+K694UFek+B/+i1ybElaKZURmQz1w0
q9Wrdncb1ELFhez+uFcr5Nwo39K2Z2eK/nmkdtbn8l/WlUoTkdwv7/JU5cf+tlCa52+1RaSe8Y7z
CW1gl5fjOmSV/2bqkIxMSaCTdrjHO6xeSX5D6WS6URmINSnmShMTfgTV3hXsJq9WkizwBkERfy+c
XlmEFcdagT1LFhzFnz8gHeg42mtwb2O0lsaGe5NzTqfOBMdTeCkzlWAYAMeA1csnKLe71Pucr3wq
OG+Q+Zar485SXmUEnKC0t2tp9WritwuaR27XlAbes/CZu9ijeuHEpucFLtkVn8t0+pwvjXC9DH/e
jTMf2KtowplBgO5ZTwqcVMnj2riucNIJOEb2a03ztgzqK4QFOQyKKK3ddHMbPNP2OXbGKEeZS7sB
J0WKmF+eHCkzKxaIsf1c7U9pBs+e5J9KAXuoDkbWYNUoC2JgDPF99tVnLq6jYBBYA/O8ixq3desH
oztFJrf+uypunyyDEi7I0ZuhaowBtIYBhJUgfX5RypQMq+QT8nmZHeIo2zqmdOXcb6MhYsb2sKGq
/KqllgdE/Fy6g7WW/0eImjcRqAV1Zgo158/Z16lr5ZUuVcZiFsbPK6p4YMQ+q+DuO78bHVk2Kwc1
PLTLliGCSQrTNZrkWxKnArlwzqMxRt7uKQus1/vpKcl61DuPqEFQT/DoIHgz2tSdHwjp1I6/UYJ0
MwhwNTizVm7Y8pTR1oSKUXm2+v2uOJHYJipbYiCxJeYvQ+74pUIVZaFs+xCcPM0hxHCb/afxm5UO
Dv4B+ngCUMYII0u/WZuwtmxVjUlySmgv5hD0e25A+Hpop4GpmZq1eMK1IgjZeIMSBDYNUvb5hvtu
V2NQDIwBJSokTablsZJieWGB8ehSRrjX8QvFxDs5ManF21zTbF95uTDhCzCWnZG/IuW7QtO6XOI9
n1qXikPJDaCSXsoX9/Y03iTzF457uSLRBpiCPLXJEgaH0EU5tr9n0NUxsRH6nmgD84TR6qVV/9oZ
mHOQQ0k5btnXv4kGdSyR22mYiifcrY/RLDuDylYHPNTqq0YarpRlCBSU3qp+RBGoVP3n+0YFexs2
9EO5ZjNkOyWvVi3BuCbxflbdmlPerdlmRvZFpvXOoatlVw8qbiQLs4TrKM5lVczRt/QQa2qauD2U
tzakKZYKq23lG5WaVLxtlf3WYh69aSCUwX24ZHy4NcFwMqKHkSUWws93bWGagGbow4B2Xe4M9lPk
Y+R5+GcAmquhXqTCW9RE/A2phpwVMZmlZgXCkWIIehYq2RKyXspIOIcHseZDeSQ9zris1sCRB6Kf
eG3wxOD8hHRPjc01/HsCkGCIRCLAvkmbtGxIlEqsOVHJTQeyU+jKiYqsf/s4ensgGZaGRhOoN2fR
jyyiQvpaM3EBAO5szIWP4TD++O+4hMDTah+wJNXD4g2Xl9hmdpB9aHn0Ta9RB+dm2suQYw4yUbTL
aFHhq08u2BG9JLhIaAaFxPuQoA4WGFx0Ck/rKQdHJaZPlGNqIQQWH/Kj9prsLNiDIzp2JDGIVE1Y
3yFYgtwhrw4ewu0kNxfhx0CdPxhtYIoiYORbn+Kxbc5WvcwlAhz0EidwxVrW5XnJKIXH1krMAB54
KIHrBL/vv/Zq2a7fw3WHL61qYvZYQQ+W1DQaNwXOUPEIK7+6WLW6NOJNfxT51S51x6vHbXI+BjQd
bazP9BCqp6L5kns1o2tCCrwEbzAvjj66XAH7NRPyX6HTsCtvRQsEXkGbefkPJe5kxPwHoW7s570j
XvNxoFA+CDTLkHwXv8cQknaMJKsGj6wxyUumoun3ckwE5FGD+QLSaVmUSurRe5yNRr8c9OCALwWj
O6OUa+yWeXPa2pjsWAVJqtH+3/x4QTtjZKM3a67aK2pE7tKPn6eMliwbs3rql/4JlF4s9wn+cOAI
z0Zdf6y/yrwf2+BeJUQ0jR87gB3nDva4DmrnaloaLIF9zn518N8FSb9dJrIC6otWHARgveM1SM8m
CEWkDHLWQTLw8tf+uz3KyF9iZcRxbwCtscIa42zYPaTE1C2pdmbXtfP5SEiKoqOEdIVefTNqgnzs
O8zIg7xYHG2wMdbq7NU2huqp75djoMIiF/PcUvY3OPZWnQ2U8KTzK8CEeeix0xxy8IptXm/TdXT3
+LKG+rsDKnEzEI4iMl1kJ4ek0qhik/wTcFrqcd6ttqqshgjsCFhe7vT8tKsc3o3tqlTDUVwm8HeV
iNOB3p/tXp1gHl98HL7/knzvCfSL/0RxYm+lWhptW2O/2ubaeTBD98CMhR2Dz5ZBYo4JJayc3o8C
IcNahoQNmIHSU/Pi6C0DU8x2OuuARSsX6PtJgtD+Gi3EKBj3SojKkqVynxqzoYY5Mjn2zqsWWva+
LkcCLMObVnFebV4/1PuCCotgZHgHVDiUrfhRjuF1eAP/0N2n6C0uGF9Qrk54ZfqLP36m8l9bcxVX
2SkfhWv/Augmi2szHapwxWDfJTOtotTwiYhmIGmDTWRmhJQIlIriD7hzwpg0mlKK2pZ2cPqMYx8B
mCsTUpxFyiSRUyF1MTJGfyXELyZ2WdDUatRd6neOmoGzS76sY2Tk18GWy0f0MLkz3ZXCV6POyB1X
+JeTqPZgjR3cRZPm/FDF14+8AHwTZPGOZkDartbUdeVN456adWxZqdecxcKmtCCE2MxRyJBwOLXX
qfB3DKfr5eQTj4y6OtJGDsmi2WnXKxsHdRwq8clo4iJH5xtII7SJomm0gF+ToqQEIaD6u7mNDTv5
Ml/BsRJhx0K8aLytgtv2Zoi6Q2jZslv5xrthumIHMXYaQQyY9VciPOB8hRYYBGA5sdwHQGOrf+J2
iHQ653KJFJz/yfwQkLWFVvt5HlFgy6Bn+oZ+HBKkSnULgBjZGOrIWYkU/D3C+6lNAm6MtaGtU8ts
ZgwR52mTDHH/FHywD+h47/Q7PPqQAD9x7DAyyBeZlShozPr713VfrPRmGbVpgFOMjwBj+rd4iMiN
qMmyDz0ZVdCGnuzUuyLoiwjZT+H0UK1glwSsQen9U5Zw9xNXAXoOXo4DszWb4h+DjwGY3LEUbiFE
5lfPVbBFo1x+CUnNuCi6AYNWekhX633VjSXSpVvP86QW0OwPqT0cGvpunl2MFnVjjmvfL4R8NZZ/
q7ZACfploF3nhzAinWYeeqmD8oC0RG5Y/OMQC3i7Alxz4uTR7IrB4W6v8+RF6dal3PcfggR83G3b
VPnlvYp5VJFfLayJjugnEk0Gh33HgkfgVpCnN092wfG5E7Fl6sBvZ7VCWoeEMpks53Piq97UyVlZ
STmpFBwgQNb1RNO9Ln7tMugfPPmT2UONJaga21ZAixIJ0L9RcyJpgyhFIQ9qSiPybtDaGvdwRJB5
W8L4036L1qwgleQkRidKV+5QxQAW1KuxXILQ7TVWHxxFKrez5wyHaMW2nnR6lzWdDyTWe4rEssET
pWLoFzxCgOiQcaai8seMyRZFwc89cJuIpWnO6/NukDufxCPQhxtrBeOrh/kHgcQGZipLC+xcZbeL
P/u8wXf4BMZJM3lu45IEnSbDBs9rFszUr9ITlf9ebr4Fcx55sEkIsMGKB3ShvgC+gn12WQfHoVh9
0dLUd9A/ajBeUdGfmGYSCp+Lhj/M8XfUTgKiH2x7CkJJAgQzppdbGEqI3ceTiqKJYqNQNa16Lpa9
spEyILcsBSvRR2WZhpV3iMn2QzWB4nJ6rLFn/zbElMJOd8HQOx+h4UjZiml4ZbUKyGEesu1A12G1
/xW4KVqnEoNCf4dPvRDhGyC9M+30NoD5knoMFZ/ZDYbs5D33o4tDDfhcTQcX3KpSsvcdVN96FRd8
PPF28l9tp52ZZg/k4k3EeB6T2UG+1O3TNNDUDaBsL1n+37eaSfvVcgNYremC6cw8mZ3NBjald+NN
H+Jl6BaIQVkdcZ4K/LmG5alsyLnItJuWuDPXb3xy3N6JnV8wg+BbcThfwkDQ+gTmYhHCoTguGqN+
9nKtrE05ZMo242esuIqrl5YRJG8XoUUdSeCJ+aKb1WVuI0N/GzdxYR512+yH3JpzOjGrHeF6fBxB
HS4WodY3bRx1w3yJSLCp7pt1Y+PrIW5JJBaq6AyXMfASK+gqi2+lvB7rbWVbuW/iWD0p4wSpbjH/
Ws67F3arHb0/pWuV+JQDilI01PZeKnAnEOa9qty1SoZ+L/NYmcVvkNJhsG6OqI/Pu2qN93PH1X3d
n/uoXzxPjHqtdjhRWsWPNh2CIOZ3NiVwYsv7vrVOzVpkEHzqWK2ojNAWwvorDXrNzjAdordaAkw2
iprwGOdVrLOOaGqqB5O1LvYn8Wpr/6ps4yki9A1Kl5k1zmYoZb5X0Wfsbb2p+VXBKd/Z/RUqJ4m6
AvYCvdPz2uRa60QsrslrUFrCXzVJVrT8QZzct2112HOoPcQWPUaTt6SJnIboC9cRwlXrjYdV6ueS
SJeEmr7K4IZbcWun3MKZvLCxU9Zd/zckxGb7ITq7R2WWKrqC58PF4KUvnLcXWVObJN02pq47BysP
MWHCJb/zFVe8hkA8uK1jvoLsCzmRjidvkj1MryxFBLUBO9aRtRJOf3Tg7OlMXBmij1jafAT5HHvR
R8qW61hqHig5pAGnMkU75dJz9KKmZm671eDxoa8/48bwLyO3GQU1hlU+tD92uhYdLd/V8OhuUni1
DznkW3P4JE/oDMTYD9uwtzIE6066MVtvWAEjgOAYhc3iN9iRkafMPnrkkU+wh2bX2CJ0czVFWrUo
6+TwxDpmAK0lnvqDaocmsfZiRS24CR8xkSDd59Ngke26MG53Ud9AJVywRKxxbSxRhJq8IyjxQLjm
JKYqooZCVsDNVPoqBFeq4pzoIHZA5azpl54ZgdyZMX0/Acf4YuoX09i+ZE6uYpSSS7bAfPzbTdET
VV+eSjMQ8ZUwlFPLiCKdLVvCF0QSxxwLQrmmXhDKPruzOmBPkPKFONNPNoN/ph9atnjAm4V1E/cK
R0TrXjYrABlMHEOWSFKaW3h4l45cjiK0OaREJyFGVLKvIveEsAuQyRAuf5V9aPr3V+E/9SumZ9UX
slu+FbrMQUKQ+0lU2oKjIU4uKnDjCT6NKADXDZ1g1xKFn3bd9lneeZ5YzFGvmG0sYvl68N0vWXO1
I9gXwqqiNg6M7tXzHeUtsrogd5RnX4NeMokCFzGqfPBEs7c0tSMyci33RRdH+S9qfL5ay0vpavYm
puF7pcxtrLf857P/LgqiABv8WRp2VtdcAwczs/XTCgmVGjgCev5KxmJhmNucXKjw77PaflMIWvjF
u3kvErlURMMX4zVxwHHEs8bvR6WYf++6HJ506YyGR9n2Ndn6LJWdpTZc7+TFaHf/8MOja5Vb65xb
Cict11Ql0MyHgHJq4uo9YG7wu7YIT2qr9NScUmkQri+VxDj29f/rAneDxYdBYukCeCqbFaidPAuU
wSdnz/1s9nG33Mptjq2hmygVXjV6BuPn+phm5+2a4WpwEsEBjyCubbAy388RW76ZhYNZCaX+zUeA
Zpw8FBaWkwkqMRUYWH8361ikVhN3D2pmdj5PD5Kze7Zww81eJzDiTpev9gv7r/8CKnR0dHFudrUC
GgbVgvsVsP10iAuWM41iYl+chdkBNB/ETrwlIHgvRyM5DpU7+WczdJIi1g2OndIwJZVU/YEN6cE1
wziFrqiyjHFDkhl00NPunYa/F+8RY88WJhZAm4G6r1dtuW9ACx9z62lQxM+M6AEkeVzzUgtRDZeW
aTWIp3Iu87uAFYJSY7gqyhqNzOzzdXmY4aTfSQARSwMeOYmIS4uFByPnautBU4lAUaa9ey2fP7f2
UNpJ3EOuFOAYSpMUlDGSMK6QwE/ar9rguZU8IrEd5XDtu/0f16J6o1F11Az/V7xTpUAVcqh+7cKx
VFG7Mq0B49YqMbIsAMK3zOzLuHbRHX59TfGpYIdPN83QDtpXb1W1v0OSfWnhvSIR+X5om4O8diFP
5FWxnmnzjBlKorEkotH7c0nMvR0hMkgZqkPxKWZsYo5VI/rZwzYLd2aK3Tzm+JZbqwfNLNAKP3xZ
WXRrvJNR2lk8l2QVE/Hvxl5NxP4m0zvQJA3OJOsmIP+eG0STFcioymHehJy3rKprH1HOOQzKUPpM
YHOhcSqMDzzPyU0pcL2BJqimppFwzuW3WOn74YlG/f60tPZzm5/HAqD3PP1fayQpdTEIQCyQODWW
Sg0/RLrwfWqkPQuuAgSvpAz5RCIJUJrpIFK5iXotnmI+oGt895VzMv4SgAug3z4FzDsFVj4jha3l
lO2ISmLiaL8GIf8E+Vv/p8++vbJdwDBJojRcdhox0IqDitmUgj8+bCSuHVBEebuqQDyP80Egu2VR
o8LnIJWzR4rNqZULfoeW+/HiQGB3lpvk4J16NPcZVf9oWH1R+bv/BjPOdGXGapTpAf3sbDMk/9lw
nRVYZsedGYYwTaFg6dgg/he9gbxMhq9irWjIck4MEpnES55M1s8c4hwIhc7S9aWvoAMngWvwcovT
Y7L4xXRh4mQSzx0LMOfch6zM9aq3JOp2W4q+9QtpzjZ3wkdKy1JLDEVANTfRIAR2lVL7yI31Rk9e
1ovBsLtH8fbJzxyqXFC2DoSHeXln5ufNBvFMufeU99/UDmi/uQo29r5rKAUXxbwvMUq8MjopWntk
Krti1ECmdxjY1vPp5O/II4mKwS6XH5wUYH5BKb/HJQFSnG++5YvQixGacrBK9YcBt1H5+ToLjkae
37ufgf8KBCsRBdQXFiCdbiN5+rArJK/SFKmscRXq79fraJHY9cTjFV/1Q3FAkUrjprjMkvJQMjN9
lDB2e30OD+APoLwoc2jksjaJP+kaVx6o/4M0t90aEvtG89kjtVN76M8jjwneqP9CE7fgxN04Kp/q
Rk4IBJrSYlXJrLJtbfjmnr6Glkzf7hb5EL77K+awmR/MRhgXxiljxPFJKGgKkijoMbJ2FulTwkHo
bIHPuY9GyNH3wUC3U6BD6LifCP/tXeKx2Ykv8zhSTsnJFJKoybPiwC4kgSblpDDxfNB/meAv7Szv
yX/iknIJllVgTPKUJVkSF5ui/uu15hzCy5UcWMtQCcj9rxbia5kuRLDoUzE5YgHyD7/eHNnbJXmm
Pv74Qu+UGHRm6mG6PADKXiNevGdOaRL0inSnFcSnCRG55iEgkZQWG2SgIqT7T/RJAj4ZRpUt13SJ
gjG2GQ2VsgwXLxnKAaUybovLoroDQMsAhcLV23D1Fv/YNSKsvxxaF0wr43ulpwG6vhSYdfvIqOWS
4NWkjlnh+rEGkF5SmoPUbIqLsDUEb0sUSd6sxHTYSi6FBf3cQoWv6UFcwk6kVBIE6bNi8PYyBvbk
Tq6HiRyS3bWe1vW+qD0JF4NP/89jJymyP0DfcTbmSX5dXTPcZXe1MG9NL3NoYBqPVQ5QcdcI2Muq
hZ0nj6Ncpldkc4AolCIhGcYouq8haA/ykVVgAp5cjqMLf3vgliFMjI9HS2rXUw8tQ0sw9GleWz98
+CXx4UGc/rXOMFfdmi6arr39dNeeTiLeBj8bxz0vVgaOIzJ6h+A/AT369jR0lga2BB73gmXWdwya
kF//4ByRELFosmxUhm+K1sXtNWFGD6fZAjgpk/xIVfCC4qDRakiP7oWDKHKKQaKtfvnijgOGQ0qe
K8hbNCayC4xkUIWdVDYgrL1qrs7qWNCQqEJCHXT1+TH1pukDaZhFj/L2GDDKbBGzwRSzKc3MJr+Z
mtjbJmMK6HIjHjABtqWvRa4G05uGcXHESYJ7EvpzxrBBUbqEDaCeNOP4eAsYOs4d2YhhUalnH9ku
mrexviHnJiLZzHSsboxW6AKjyjCBujmCYq2BsVaDdc/AIjn8ZysIlbB1GA4ahqD/DJ/ByyQcbhbZ
Rp+nonXAKfLXxRRlY2cxJWwPDwSj/n0dg9WOdgKllg3HZ2Nstre6V0MF7iTSkZB/pqfF8Piw7QVg
95fjols5difzTQF+RyHF6h/oSW4iM4TEkgWLQNpBgAjgBHs/fUN7+Y5m88bpIl2uQ4iRSK2CRFnM
W/qhWqbB58kn+BkRUwGK98yLMgrjr43K12Y/1SpqLMI2zY9O/tP5nU7c3bLXPksXWwWIZjqjEmr+
pr8Jvn0LK0S0jBiwXa3YKk/coK0S+T8PeUqJiyJCdnLxbJUHNyvU3QpGXrsKBwBvBWTYaxzcVd2V
uUwAfn5yTQdrQ+NNMqypcfDXQzE4nn7JvSz9zMgzUEVdoELq+Qzr9GcyIsYpgy8hUkbsUF3vPQ43
n4yeiXWL/um8Om12x+Bu8J1hYku/yrmuagXwf7qgNNprppegsb3YrsUsu6s/kiEtKq19YpjM7Mnd
WVNa3eG27bIYQEwk9VKcy07q1DjpR2hBcl+5GgDGRjjPo+Pl+KNmaW8/p5PqbozWouQE0lrMK+rz
zm79pxi4aLK1xbMfLLYJJ5vsEo/V0qC9jl8hUBfn/vaSjpqaRIh+e2w3ZFaQRbkXo+5hqa93vheO
d70hXBw0vc00hu4l+ouqRunU0gomJwExTs/YYFXhTe9mlUMNEHOkroh9tKYyPeDHPmfjPm5RE7lI
G3zsIZmb5uPLaTZcAOeR/kY/UP7HqQg+sT3UUcl/jXs8ZVbE53KemafkkErvcH5salxs+m5usFjT
LwWGWnawe/rJ3z3n2OlNQdbXagpmz0BRlbfpoWmQf/aN6VxRnHvLXaRzj2vnwYdGee+AyNHVREpS
fSldPdv1ubUdZAwxYAREu2Rld3zrzDWJ6M4KNp1NT6JYM6Epdi+lrn5oJE+QTAVymZCtezDqopH7
SpaKLiLeH+c3xhAExhB+ATERwYgsUeQxDe31YIzqkeY84yqPTBeLryBnxBYL7I+vza6ubEaCLc3S
zfLQd07F5Whk1YKHlKzR9uy1WOGsPOC2d7HsfgL+I9ovjy+VOsDp7vQc4rj/9yWsBlncJvLrs3CF
mcOdyb59HJRsAlnpF7+/axBO4FXtjaCw1Wnt2sq7EYTFZALRumPaIXuDlwBSLj2Vitt4lR4U7LE2
TNYpvjIsjBacVSFE8nE3V/vTF5Y9b9HaGtjrgLZznYoFEm8ypjVU2KS2TyIg2hiakz6roZhGaHYs
bCnqR0yQKih5MloDSfbhH2yBz8gnTyp/3OlZeYykzgwkknaENQKoZOmESoF9pTZaIV5yRc/FogS6
bj9OrMwRS53MQAORk3HbfwPZ29WZmWU1Ma+4ue7ilrtWAuzL9NFSkBIhpOXoSSibeuyXk848hX0D
bnrbxOuK6UpNgIa9iCLtQBq/qhoGQlEPNFyfhFDMQras1gjfqXC9PsCW5uQRp139B5DILVQCa2IP
L0cNePVQrdMNl4/SZS1xy2/li1jROmZVaQrGcXYrjw6UCyhiorVhw1AX419N8svC7DQjfq/8YHDq
LkFsgEXcGc+6RkhFUK6pv3NovV/EScImA7Cx9RBTbYkv3ciIglFjuKlQ0vy2UdAFRVxFrXjJGRIa
eVecetaZ7yGr25eM9pQtkke4o5KQczpZTOq/9SPhRfqzoLSqPKTeucavBCuqOtwO5//mYw2GWM6C
6YelWXiEUcaPXvbDpOoHqNaiPG+IrfizG2TNaRgT/tvt+4XKJtWouI/MbQ6Ec5LOqeXXEGMK0OqF
enNCAMGaP12C1pWuu94nF1rk/ai8jW6d3CGc/ZeIuI5ILAG0V7KBJjgVGDmtVSvMbvCeQop56BdD
NvebrWda5BxiRme1sYUYHb+aa/77clALw0Cr6VbSSzXTszJ6GcSfh75j48Pr21VuQCw8zc25UH6I
qVsD0F6PkWmxd/o1atOXLhSsOUCEg40ZpxqqslVmdxQ9kb3ytEx3sV7eRwbhT3J45Bjek0gdJbcc
sq4G8o+zGWne/z/jtcG/P9peNuNa1gt96B5fUQDs9K+7Ix9aTaaALaT7bAqAidaiFFKiyD9v0k7R
9Kqhp3ElDdDM0GpUnva6rL5as6Yzo4o3O+krR+SyhDbbR4edAdsfDcuza2Fbp+cj2Llp2x0iu6BS
9A3nqKmEQRF7Z2bD0AqnWEEoZxRoWFPQKR0ECmKCIlBgJf3ZUEQYIFJp96vHfmy9dvXP3xTJ8H75
SrwbUa1xvmWKp0q6mUySwHMTTKJ1fp3Nsk7EgPMW1VP4vJmIkVQkyZUEWjmjHzgABtk5EHMVgKOk
0kLCKFtvYf9V/rlY+x67eDpwFZ1NDgNncEkYY7mnPyzWIV36AwMtgt7e5SY69qmjava75/h3BM9+
cD2RXK6gkl/P8jtQoUGgMBGzOCYHXJRdIQJquZeuolSSG7pvyvl+xQfjHbO+yjQUAPsKWR4LpxkS
a4mheguH9r3jOhcI+oVPDbgTSudDw1xBKx8frDwwuw1s/U8WyUm+qaXFfEgJ3EdKSUvT3/7L2dxX
RKIDkQ5/k0l60tlMno04zLOVJAGoclwqaNdC7XbmbLgBfl0c0fxpq2GoIkShQzrC6IipZgWdbydH
LC2f3TRXAFAeSDmfRES5RRcWPGM0uj6tlDl+8YCsEDxcUAwFhipJAyd3awtgNOaE1DTnJ/FrRwG7
bQ8spELhDLtw83lgjqPzl0ZZs1HvRiNjKwBFdryWH+w+mfQcJuqdkrg9Va89smualE+5BkljDG4j
vPMc8AbNAOaSOpvZTDrC3nyIbI7ALAEFvGIRDcTMKgKxCS+rabaTz9RfFTXxoraNf5MfZQSDavUT
5/EXoMImnh8l8/6TXaKBB9Ytzi7Au9aPnpB8mwRQXcQVeq2MwRR2sAzEQQOYaG8Amf9+3MNlfQBH
jGuNvk/oimsX9BU/SNp53KFJvrRIdvPaEuIgjQCKhfyS47ZwGRD/mnlOTYv2EYayz2PpQXafq3WE
fd4s8K/ONQJF8KyLGmtEzjuYSFxHoEBEOD2FsEJGyQTN8yjt71NS5Iadf9zDlNKPrsGh5KLwGs5p
5jDPfOTe+JAdgY6KSgVFVbCWzNIBoYhLz2ryQPZB1Fpr5wyeGcxMmazrYqGSo6gXzn7kNsyFGN20
arjHEXj8wHIJC1IAafTjNZpHNPSDvveffnltTzAZTJaIVo03YQ5AqbeQl1l4MiIdudGmV7ua1Qrq
j6aAJId0FtSsdA/v+WC/Ml4wserkl48QRCbBOipksCIDHLJlSzsPr+xg6ot2ZFrM9c5o1efhZU1w
u8dbZZk3NFJrzf82mL92wN/EhjjHyW01RhqzRSNZVXi4DGp0jk6O1YwLKU5ysLP1PANiyDET1hFE
XsmQOdlfESR3LNEsRYuFuiUJAuRz/038b08n755c4vegMlXYOS5WFPCye9snkneec/1aADoYnFpb
praHGKbtAzyoFX5/Dm9oXqknq58rigTrmZceWf/ZFTs30Rn0ZeO7IFQri2YMk4d6YpLQdiydb5F+
kScYGQiE7PgRkeeheJLUgGxX6oVpuPdMdjY/roWJiIJzUynUN1EJpwaZkaF6skS9A/KPjD8a97xB
jVceznNH67HvaSHfacXbLTynyAXwudY4CB30SL+QQv0Ghw3CDfFiJhwfApzmp90NPPggC2w9Mv+j
KxGLDCwMf8lUtA4HDtmN0u0qua1gJ0eKJ6Ur2w4gXAKiMKskd7UzSQeBCEAdWvNNOV6qtsqQns1Y
oGlH+7lHUe0gjKjJZwnl6RLPZ7AezNX+3+BUdmm+sKqLj4uTJ6yVpiA+FzL7JOkw9iyHGzQQCMyD
bDR6L75/ZPM1qcyBNs5LY9ss9xWJ2iIZPFedMWTgQJJqmM7zmpj7tGftboS8od12z9c008d6fWE/
GNfuRT2OCdDuw9fctlKpgil87NyUMFeHwHj4AYPlS5ACA5Rh+gVE0BmKrVcbVZ5jxbLT562TvZ1s
E0om0KuLh6DhTbVRm8VeWWuJ/OydYoseSaCA/3dASnT9j+o9ndRVKXVUHrI3OzGAFcnw2q4sCWQH
h4UltwXjndsu+n+vPv0T4DOuI+MgTU/PR3KEDDYbvDEDzQGYQii0jODWRkd4T190OJ5oS2tOOGDE
xvEsAmJWsrbuCNRpx69/r2sNnYPQmYmdso5neUk+CBM6OYMdUYZzpKH8ISseXSzecXrDPumY+M9V
7pnxuLPTMgK2d8eyrsXC6t6qSokg7IypN+T00x1xMz0VDPEo+XOxbfYsR2XrnI5BwUA8QwD+aRit
7S1zJzYXVxf0nEZkFkCMG/09sESWF1hivo4kf4sN+zXTSnR6g5xqIGT0nD+1Q3UrYQgmADPa+XN9
H6h+4VtXQhEIyjml0J+MUxq2Q9H2ZcAy0PmghV+6l5HZY0fsqAh5pNXoDY1TVQTat8xh6rZc5O/G
oYd402QSF3u8tu8Efrr5s8EFDZAcAuiDLWXYyTBLGz9LsYKX5xsxzo4GPrKFjWBoDQt84KAsfzkP
Y5ugs6KZGXeFVgRz5TmeFBOLLZnWkRT2fb6CwVJp8JFuYU0rl6HlPLRou/mflH2SnQsplxu6irCW
Db/9NEkG9HFjk35KYg4QOoQ8LNoUSRks5BhS33ZddUAGtHAkcRfMdM4ZoMAEn84aUcUDr5Cd/T7g
2KziuF2ebSyB10TkzR0j/GxtTiaYkQUB4X4ac/RUNlrSI+a3YsmbWaFt2dwaannW0uPmaFCK72wN
tu6Je3z4jxI1Bk0p/QFn7KXw86g636Uxk1MrZlCMOyH6j2ZY/qKDd4wlH6BqhrzaidKpnmVZ1L/R
0nz8GQwOFgiHITwOi6XDiAVesCIFBpve/1ko7WFEa3F33zEHRx18Mh96ttR6DtWo9LgcmnA9tXbo
HJI+oBDY2I8nKZraa7jeOYNi0CXRiADoVp1r5eDpE38ls/8rhB04Wi7/AuqsLBGHsh3QFP/sWiwv
O9RM4cGLO4myLIyYtrvFTxArif60T9ALYgHz5vIIN+lloANmoQzC1oW6Q4T0vEQ3cKtqrgV/lZdg
9pj4DFoqtwHMsNjbT70Hk0/lektk3ssiHyOHf7frHeQQpt7Kr7oB9QyNEMvPy7pzvZiwXICKjGuR
BQLVOMRtU4Ocps7vEBB3eK0zDmjbnB8cTihQO1HbNZgDT2lbKM3gyBurR9PXXEGwY1X3FsA1xa8Z
dAnxQBJpoCP0iunOfK/dAinPQ7TnR24F3BkKUFVBuon0B0+414eUHzmlbGaIVL1+Gbd3PRM62z/j
iP7l+hqWhbrGeQb77quF9rxBi5Ux1nVUjEoNjUfGpRbXGv+PP7pDXdH9PTlGGt0aLtDeH70mfWFy
QpPMnlDG06MPWQEzkz9GS8Gvu0Hlv4GAx5TobWgXlZFNP1Jtinwy1JH+FtBoDaMsyTdqMbLKrOhd
AKUfklW84sK52FhK7HZJWn83D+TBH67caKNMhuCHqX779Lu+RXvyD4hBrwALuGJ3CutG8S0CmEDi
0ed1z+dOZrPMBCB8WZJKMpuHRMjbLP8kf5cAUY9dLEh221yIDWuV/ZbwaMgYxbchRju6f6M1iqdI
DGbEjzfqI3/4mHO5GpN05MEpAAFirVYTEoJwIQKV5JJN+8UdXKaG8Wt5hIjya7VPo3YO6AUFE0r6
it7QGYQfQDRwEQpU7nVZyfvoGqm72NHjC0Gqrz01CZ3Qh5q+mSQculwFGhfqmqur1up9jVt1rGz3
tDkv3M3Od+LwokU+Pjl1dxcz4RxFLWLeAUbM0y1S/BXi/xlINP0lyL91/NraTGZWo/8EASbu/G/Y
1VNyJ4vWig3HUUhU9q2v5EJQNKUsjsAnA3PNDLLNu7HESliQKjRlRv7b35Na+ySJkmBHpVGXQ9fe
4cwMdayIyHIHec0OFuuxlj2yR2Uzv3ODctOtAb2CPL6TGJQjt86WJE4ZowEvsO4DmolnYgbI9O2I
lf5BvpnbsfJ8iVJwtlmF+4zW0oqbvh+af1aVbdHDzW6PT1bsI75NmXE+JAPytTyUUlBMTUnDCf8O
w/IxHIcKNpxc/ylzogvRYtHKeDKJli6Dsbf67F+34N/Hqu8ogU+EgbHDIf2IWFo9ZV6SgCB0KsUo
kqNjKRCvSE9gY69Fj4GBPKqOjNfDoM1WkAbGH1ruAzxmOBiV0ZWGtyLkx6yq9FvkKH9pxsCHBtZY
M8NI/1aUCLvbo3FbAVfS244ohf3X3hJnRcVL0VjiU6cex+qy8aKPmH+LUf49cAY8LYgf7plIUfaj
ok6/6TzJMRhPuJrUYFlopR1HCIyaLMoruA+MQTt7oN9Wkht479N8AI5t7WF46ci9lw8L847W5WyY
866EM0RVr/ZhCMASnd/2rEqeXkxYWRR6JfP2kOCLsOu5B+M041n2+2ROEa2EoR9IUOfTpWpVlW/J
eVhz1nLBVryhah33HCWAqMLsK0TlCNC+B8SVCbQ2nGN1vU/LQZzkBFQjAv8Si5tC8iopfWcyICVs
gain3GzBeFCF+prV0WmEC9lELpwf+uD8vpACZg9xKE40jM1ew+DJAuBrHOj14C37YTFFnHGsRoOv
35N722UA9F0UbwfmdePUMb1i9qr0kRxU0agl6CpIGMHiS6dvPcCDEE21Cv4TyHVz4gjeW9quIXTo
ZtOR6EpBGGy1wNj0JE2YGKLw2/pz9odmiSVTOaTD82cvPMxCLRJNBgBHjhv7AFF14mPLBUKVjyJW
rwplBW3ejvGUHRXnIIk72n/QrmeixcvWOvFYrZvOUOCBEFx511JkhyO1ge6iJOUPOFlRcSgctuss
X5PgKHYMYbp0mEh3AGiqZc4laoBZ9lW+Xr6dAfrfB+gRuyTzP/01P5eb2Po1m6DKL5aqdAOrCGMt
+0oqefgPoMLjpGy7aNsH/d+cr57+A3FimPyV6kQjt40Re9P+HeAgoGSDuYhuycNXOGaJ0d8WPTJz
GN6jHE3wdvlnFhDRhu+SVZBbfvxqp6AAtViOoNU+YydZ46xUxkQX37mUsKpQcDvDSof2yRxwI5KF
zLjnNJBz/dM/M8L0RXd+Dop+9O/N6TyEAktSXJqlTdzmtggLzW4x+UuYnHff8IINF1yO05dUTQGx
pVnFGoUM96V9I98Jr1IxQ8OU4pGwmU7InFMPftWcxKCWQBwjV9O6vmy6LLA98nqbksB5ViaXDFb2
y5XvlSwaSsqU0/FecKSKYhss25b2BcYWGfx0qryFQmL1vDQnO2gu/LnLAQhyxtvGGmUR/+s+cTEV
235IN/YLozFSN5SorYv91DCv8dZAPZGkEiA+M3dg+K5XEFlmtsK3HiadaFJATVoJzIJFnFtGDPoS
z1JI68YnO8Lc3g0L7nWdfA==
`pragma protect end_protected
