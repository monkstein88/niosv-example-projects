��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a���5�_�o�73��V�i�EY�E<\ţ��i���ќ�{Y��v[3H�=�"�d�.]�v��+9	�~g��f&z3>�~��̧:od�<7�U���Ѝ)�p��h1i���"55a������۸��4S4�>q�&;Zd�3��*�5˭Tڙ+?@<�t�S!��NZ�,�F=UTLe/bN���F��&�,�7��V刻�?�;gj���摼�kO3�fV���oH@K<I'����n{^*9���!|R��K)s�N�s0�aI�0�nR���c�@�>¸ax'}j��
�x/��}����7915�q�
Vs�q�43�֥[>�G�:���8ƞq^�y��:R���D��Ų���+�b���W¡��}��j�KB��E�q2;d���qr���?���<�n6�Uc%�-�O���Y�8g�P񶭹:��0>#WW1[��m	P3$f�Tk��/5��m�r��i$4JW)��}M,f�)t�����ۅ)~�C'��R��Ig
�����yٖ� �Q,~BY%�6�6G�
-X�д�8��%�\_<�p%
��]6�X`0G٪ozĞ%)f�Z}&��#�����
~sA��T��`$��/�����1π]S����:u�|��<�������t��j��QW�[Y�/��D��(�|������7����D@��'Q��R�j�d�J
�D�q�hz��)*����Dv�/)գ�W��S<����}b�~�/��z�5r��!�H����}��Jia�.���BhK^h�����-�әㅮ�
�p�lt��i�>�g�M^�^-)N�j���f���NS��0��2F�z��%����f�p���{�e��e�B�C�Iȥ�f{'ę���u�c�Xp PԮdOIߊ���U�U��Z����`�+�cIɣ(1��$�2�#�u0��5X���&ZX5�
4����_�� ��R���V|<P�2�W�MqI��Ή�[�1�>��h�F���g��(�(�5ܦ�;CC~q���Z&��xX�،���Ow��A����k$�.���o��>�����Q�jZ��!�@-��y�]�"����tr�{��s>7(-������%�]Q��׭3f���x��7�@̆ʚ��.��x\%_�G�h�Hc�`��%Z{�V�M-�? �p��a�~-v���0f���8dh�Ml}X{��Kq�s%���ޤc���(z�C\5N�F<;	�����e��}�S�@�*��+�����2��o��H���V�jѝ�m��@�rAZlC���F6������<b���!���n�kڷ�8g2�)�8� 9����v�6]!��k��nT'�v�UBx�i���x��ٍ�6���+&˟��	CfI���S��D5F�l�,{2u{;�:��*)k湱�e3��sl�I�YZ�+<�\�Tl�glK�	�|��q?�
�e1�#�o̵c�բF��a�Ɇ�]���0,
��q�pT(��M��A�0���O^%jw��d���1�r�������睬����佅����<)�	,Q���\\��vO�K�������K�9N��,��t�*O4TS�a�X�Y�}r��ߐA��f�������kw=;x�:ݯ���υ0�m�����΋�~�;����
���B�|�ʈ��b�I��q`��A�,.�Z��'��s��I,?����`�|
hl	Z1�j!5�ZHy�YQ�刜'vE*&�X��S��g0B_���QjgsV2��s+�1�{�+�}�_~�'��]�&ggl�P%9��������ƃ��p�ZtM�Ql�M&�� ڃQe#�cl�� �����˽{B�ԈvH���� l�snK�}}�ï�G'�r�X�����R}}�r�8/S�:I?����1����ZQk�gu��F�1eW�#	��d�btY�VI��猖W�˔��$rT�l����t�B�M���aQ�m揶	Z����v^���H���جm[�b�"�<rE�y��'>�6��z]n����h�N����-�K*1>-k]��ʐ�\��g�'����ğV$��K&��m���td4��7��n�0>BT5�$B���`�.����'�L��ȭ�?�l���N��}��\��P��)ި2�e�m#4���m�E쿕.O�<� ܍5����q[��>�\K1v�fp/��yr﵄�zf^.�Z�QP�O�|T�S�DTOwʶ9������u	���J]����*W�������C�~��&k�Qc���E�̾bc��?�sT�2pߦ&jw����O�c;�H�S���؊���I�j�>�?��yv·v��x{�� KD/����?{�z�*�w�09�����dI�l�w�t5{%n52t�ю;;�}��9��RQ}O��B0tؐ�"�yhu����W�^C�U'w��C���w�P`��{T0K�˘��O1-���1�dh&=�:��N��tǔP���b7��}M�yr4��A=RL�8�8�#�O�Yo|�=��Cb�B�-��M�kW�\r��lA��"H���3��?�,@�ߒ����k*�1.�$���_�:�����u�K�e,��]� ��{ ���D��G�'�&����{���q ;�y��
W3����]���_�oa�KCU�����R�&o!��WS�	=h���!���"�K|�	�� ��s���!H��"=�
��vQ�n{WpZ���p���JQ �N����[tQ��ȇ����:D˰��Z��i�p/D���"G�	x�N��z ��EC��~ڌȻ�
��������UP�)�Bn�el~�~V�"�����D(��t�vq������ũ8�Sߖ�诊�l�n󠓆YF�bX�1P�f��|�	&�?�3�I����~���s
�J��2{�5��u�$�s��N�ȍ4O?.��|M!�7�g���R�%D��]0c���d���#Z�K�la5��,2]9�H�<���ɖ��t��ӏn��\���z	��' i��3x
���g�����e`���bR{�A6'��9T dUy���3����g%������R&��\l�c�"�ȁG`��[~G<	Ld�3��z��C�Ɣ(rوSY��{YX�)�^+�0�j��x�|��G�5�VL�$ef�R��#s؇rPtO+t������&�lʐ[�Q�u�'�
D])�b���+qY\�]��� ��PRX��"?>5��y�:��ϴ,6V�4� ����H�%,���m�ƣЇ��cY��DF�@~;g������nӈ���)U~����ۊ�7�0�[��$�aeq�jW(]��?�{�C+�Ed�0�6&�6����^�7�!?N�-��ָ[��S�d� �:���P����pe��j,kYEe-�/<w���O�Jp�E�˨�)$���; �($�s��"�&�n���P>�7��q��~����?}O���'e���9ƽ��!�.�6���B�o�m�3�����s���2����T�����^��}9Lp�-]�ͩț���m�Rm0*��P��ʄ��B ,���ծ���e�3Pe(:�|	����I�+�E�,mKYm�`}]�bU�O�����=�OQ���Ȝ���u�wpxF�B��(�^�8��~y��wB@�I�M�-��l FH;:�W�}up�y�i�/�Ϻڜ��1�y^lp��~I�}@-,@�N�"����}�q�G��w7ļ�����z����s$�SY{�ɗeb�,��d|���!�hqZZ ף�t�����ǿw�i��������a����S�0dr�С$�g_�~�|H	nshA��Հb�hՎՕ0Ϟ����(�̕�VS�&�'���t����SW2?��,>@@�D�R�k0���ϕyyҝ�}�.a��ƞ�8m�y!�<,��Ru`�"���	��P���<i���௅ڶ%���Z뵯�L�7x��j�8(�2�<�� z�(3%�?9��]�����$҇zA�J�t(-�
��_�g]Ԝr�ht.�>�]�S3a�y�S�[';Oş�������)'ON;0&!ND_��wza"�򽥭���� %��n�S��7jj������$��3���X��@J�2���%l�ƕ-�È��QNF�������}�/�I�1�3v�����Cݢ²��{U���+�5/�jLX�3��il��S�R�}���M$���$��T[=$��,7�-"�ֱC��L��A4�b���~�R+庱^���Vu���S�����Q#Չ�^�;n �X��v��j+2�GqJ׋��Ij�yNN�Y�j�e��#; �AA�y�jɑU��W�9�"�#B�S�Dq�A>_ˈR��u)h�dy�Lm�2O��~KFĞ�xGq��aZ��Xeq?�Xf��O&|<� |��S�a��>�J��i)���3���~�q��?�.��Nb����H�϶[!$S���x�p?�0�67��T?5����ܙ�lt��GD��]�·A`����kOR���
�5�4��(��Jʙ���V��N��_�0D�D}�"�@6�K���pfEE.�,AU�[����pƧ���U���Ʈ�=>��غ~If�Փ�Z�3��i�{o���� �hv����g�N��Rks�x�e����*�"�G淨�2N<s���ȱԈ��ҹW�tCJ�`[�^�������Hxͦ��>�4�wl��α���1 AR���3�t����H�i���k*��ۢ��s�eB��H'�&wp_i7���}���v�����V��M!`������lz�M
m����5�lsO�&����;��#��B����_���ұ�4�u%X��U�za�
\����!)Ѡ����T�d��N�U�|&���Z.r�`q�G\��.�Y���2l����Y�ۢo?�4l"�K��1�K{��˟�|%-�T4��I�ܹ�YI�}k�A�	U��m���շ��+�HNTWmz=^w�������@�6�W�D�����gg%�)����9!��\��¾5����OU�I��Ș���F��!ꋔ��@�of�ь�}�q��ħ?���Zi���\~h�3�1�)o�*�Z�/�,U93K������d�6D��8�x�T��?�e�y<��V�$�n�!.L&@�aANp@Q�<t��������@�B�l1�p�Թ�S��<��>��]�T��
<�e���v�e,�i'���}�q��3Ξ�M!3:hd7V��7\.F�h�����T�Ue��,�~gOy������y����_��$a�D��q�shi�!0�:3�2+t����)���e��."���50An_vO��lW� ���j�l�j��G7�-��+�4
��5C��.��-W�� 9$�����<-h:���<%@�;J�8v3Oco��a	�����6�}|dKq7��=�L���S�5��x���*�+e���@Õ�C�b�5U�8G�rHQ��Cc&�F>���{䦟�9I&�i$��;��6:Ĺ~R���ΐv�f�GP�u�G�x���1�5��������<dA�h�{볍[����r���>�V�~��A���vd����lP�,��	�$A����Q�8�؋U�|��\�f�sʷ��0���~��2J�}̤W��"�M�����۲����0w��B��cV�x���[bn@�)�ۈ|g� ��3p��5��ɕdX)>��)k��������4$�˞����Q���Ŷ!�	�)����.��o�c�Kb,���Jy�p]�\��c[b߇K@�]����4���ch�,՘ç��ej�Y�9�(�o��=U��9�����ٙ#DH:4]���I�k��~C6S�ɂ�����i]ցf�_�΍,X�����k�i�{��KgO^�ZS���^0m��p�q�n׃�w\�=�e����!�S=��ƃ��B�ޱ Ţ<�.;\�jZ`�.M�g��l��� �r�|ǜU���4q4T�-K��U�r� t����d��S�7�9�^^��i��s��KcT��].q�N��ٷ��'4�(h��?5o�v�zh��.�-�~�FM��i�m�$�=� ZV.���͂����0<K+͈��u�l޳��L�Qv<�MÈ�v���H��e1��TM٣�$��U�PR �%�����
�؊�J�R\N���L������6�.�G�M|�RH-�S�50H	��U�o���HmF��|ѣl��H5��Oc�dLQ*�p��.W� �#��#	ew_�d�W���r��Ũ�+^�j~C���˽��\�H�OO�S'_"N��
|(���C�|��Kߵ�F�aG�`��DčZyR`NB��-?���s��`�WJeT0�WR+k ������t��V���q�T6��f�܉��_V�9`��ug�XM-o#�{Ĕ�����})��s��[�e���go��`�i�HTu�dS�eE�kH���p�lExP�o�
־����@հR�E���[�x�!׾��B=��XfEA��_�n5\�\�U�Of0ClW���[�` <X۾)�H�(ǐ�wB(�9��ںv��Ǆ���`8���4&7N�����$��j>�O�z�t=݄�9ǋ�睡ڃ	ʭ���k"���0��NO��,��[�L�(��k[�!�@��x�V��_��Hh>,P��\v)��	�E-6u�P���p��V�f���C�p@ �̛b<���Doi�N���Bɯ�Z<4�{2`sx��}���R��p �+�-�|Y#K�B��3�d1�qQQf���վ�I�[ݍ(�����WM��8�PS/�.r9Dҗ���=�������O~ຂk��n(��W��(�l�<}�K�_�hJm�ԡ�9��yTVL�Y�n!PMo%��#���ټ�4(�޷��tK��3�s��lKfo`h�B��gB�^!
<vr���O�`#>�+`�E��V�����h|�MP�Pf�]�|��jzm��z)����A)T�)m ~4����+�xڌ��cC���En��"C�(Q��Q�p)n�O!����U��p���k�<�\J�7�Щ��v<����!l�>~P>�n�\�l6Y������F�)�_F�Wͭ���%�[	�lL�)�8��)��.�LVWWn��o�W�^/���+�ԐA���$Ѝ�ٸ��/6\'{��Ҩ2兴eۙk�e��N]�_w������ަh���RE�(�O%�Cb!��Ch�J�;^�a�7�ef��m����+�$CBW��+ݰj�ymp��M�2yD�M�T3�2�z�6.���̹���`_Qz����:A�S�	�y0~Ҕa̷^I����-V8~���qI�$�9��<��N��Xb�T)2�����%
9�#�lC�B��@������N~��ܧ`�������"Gz�)�|�#e���-�{D�%,3ym�ˠ�E�����R�.��I^�?sqU��MUl@OޞK�X�"�̱�]��H��ޟh_r���D!.�{��t�������S
��d�p��ޑ�� �-2��t����������t^�ҘG��q6[3�R
I���O�k�� +�j������ 	��=`G�'Ы.N0N��#HR�(#Q��~������z`s�2�e�[)L6ǃ��`C�H�9�A�3� ���z��w����U�q��������b��)(��N0u�h�mӆ�$�;��\
n��/4 =��X��°L	X1����:�T=���^�)��8��κu���	)=�4)/�$�8>���>��@7�J��5��hkiOf��'@���MmU�ڍ��Z�b��QM�鐾�K�\@
_~ۮέOa�G�r ��V��o6�5�AAP'	0磇rJI����Sσ�-���Oh�<�_�$�c
���>�)�Ő�Ȏ�"�q8h$�d�?�?�D�;�d��boF��T_�@�#"?%��q.��d��Kx�G�2'<� G=�z�H�oCcr��m�]��zO9�%ܙf��m�"���6��ź�u�T�_����ɥ�#b�� ��2�� �T7��%�b��=�3��3�9#������0y�2��?�����PE��$@�#��4��z��m�W�B���/f:��T��+Ů��ZG>���d>�m?���ׯ$�������s�L�;�[�D�.���4�'ݪ��� ⠟�C����� ;�Z1f����R�k5�#k"?O�0��n5Vj!U�v��aJ����xmf��CRG�E��u�MGR2J����`�?M��猵�aEr�@R�ӌ��bg��6��j��h��潆������tf��J��a-�j�i�=t��\��ټզ�|�OCFj��gj�kF����2��e�pj���M��m!�7Q�;8������������Z �,I�"߻X�xs6L�"9a�}Aj����nϠ���F0:L��2�
I=��ji�@�\�g�Ef`o	s�)�sGi,]f��4����F�/Ѩ�'� -b����w3�5?���O����������
n��\���;���.W��I�헠�p=֩y��]�ZM	y��t�t����~y���+���A���U��w��Yb�����d �]֕J%�n�� �D=II��T��+ꀧ��?�4��B.R�r���/�3saZ"�5�G$�kb �1�����@<�&��!��Fu|n�&���̽�IRh�����9~�������5&&V7�w��VCڗY`ࠐ~	ҧ����Uz�ɸ�����1G����	�MEZ���+�7��n�}C)�Yث7q7�	1�
�@��Pl	5���Ө���g0�Р'��3(�<�N�𩔝�	[�<�,��u��ʧᐗ<�O����5����p�q���T���ܖ��z_=���^(M��!���$��"k%o�8��B΂��e���'�E�x�gRՅ�h�W����,Nr��,�qV-��Ӫ��!\��eűv��)��q��+@	��=�7˼�7~�,4��0F3�2=��- �l�C� �W�Q9���2��W�`�.\�6_���`��qV�Ӹ��A��]T����$PE��I��p�(��5|���t�i!���ک9�ԫؓ����������p�� [{m��<3��E���-6HU��O�l#��z7mU~��S]�G��A��i4��C����7�eoj���c�|�Z<��zw���fP۶ �~�٠R۰�1�G o܀�� �H���Qh?����U(>� ���������b�u��^6���ClL�e��z��e���P�/�L�N�tU[D���q��`�\�*�0�Y �����*���$����� ������J�ҩ�w\�J0��q�$�M��V��ƕ��. ^Å����g%>YN��� x���J�3$��2���E�x�3�tʲ:���������Zz���w;[�(��<'}�
��w<�Bmu�??f�3��ì�m���oR�g"V�M<�a��91%�7�����j�9�߸IK,����$��I���O˴'����N\���r�"��H�4���5>W)�2F�����o�WRK��c��7Q�m���1
���[��.l��(� �^%I�e���e^��>���'q�1U�A��.}v�)���½4��a��8l��c}�X�������?��C�*xdfX�f<�:w�����(�_J��ҟ�CaH_�����z#��)#.q�R�t�@q�[i�J�&+֠W���ŋQe��J�h�(��oe�Ű��M�#z�P���E{�j�����q�����j����֚	*���*3��-�r5��&�#�K�&?����C?���#oI�e&�Hqa�Ntx�v�{1�}ж!"��m�~�X�EC����w��@���*���Ǒ����u,�˥ciS��	_O0����k�(L������K��6#��3[3�;�Q�x������ﯶ�;�� �0�s�7l����hwpј�tHᑝB��c7�ۢ��Y1l��M0�8�v�j���d<S�{!��`��#�阼�����R��Z�!h�����9��_\X+s��M�E���$ <�?���"��1T�[)��}���EG�0��/!]�B	� Ɯ���<}).��qvA��xPt�'v�.$�LA�WF������0� *n4�%#0fpYB�κl�`0�U�p/���">:��14e��ζb77@�A��W\�;9i���>�F�|#��`'�d�G����'MZC��H�E�1M�NJ�h�?HPܢh���H�0Z?�����r�kD{���`�x>�ٙ�+6gAܺ��.8���=����,��JQ���L�-���R�	kd#r�����R�1B2�y���%NiI�n�n*��՘����+�6��|guq�Oa
 �e0�� X�K���H�|�1?�B�Xe(bB٨�R�	3�#�XC{��4�Œ���5�������l��b'�������r3O��_v�*5 5���c���/g�p���������	K�q�\�yKg�
cc��Čc��
��<y�S�|}gKwS*�L����ȍ�A0EW�9�m����6̕PKԌ�V� ����K0�l���~�D���*�J��s�|�pf�N��m�%�j��b�� T��~�ܾ���R��UEC��](P�t6gL� � 5x
m��Y�W�`�6�ߠ�r��n5���rU�yb��B}>�a8�	|�c�}N��S ���V2nG��5��g�m�4| �Ø�N�&��t��TXx"�n�WQ?�� �)Cl7czoc�8bO�nU���;T^re�_=�� �+%�R_= z/���m�\����F����q-z�`E'�.}�U4i@�q&�>L����}�ڝ�<��r*E^Y32�]�"5"�T��.���'r8<?�^A�Ȱ2�*vWM]��N{-3y�}��t�쨇�r�H���`8P�(	[�&&Z��#���`P�z�1#�ǋѡç�q�1��}ܜ��s�~�b�]���8 ��厹>���qķcPXZ�.��9]s3�s��o�x��[XÅ�$���]ǡ���k��3���>J��R�hYX��{�0�уf�SgV�ԏ���(���'MŊ�B�x�J7�j�:N��gjctv��PL� �_aҖ!<�1������":���z͖�&�H*��P��2�(��\fx�O������r���\����+����&
��b�dܯ,�7�l�s�K>��h	�'�R6���ծw>�u���G�:�%c)����xu]��e�ذQޝ�-a�+4_�]���S��H�uL4n	\�����k���Rt��=�} 2B��/z�Cr�c�3�>���ǿ;t�����._��]0���b�����C��d�`���`j��Ӛ]+0�#
Ԩ���f
�Ԋ�˻%��{�ԍ���M�'�0�8�׵��	�T�@��3+zn��&v�/��=��i� Y�����(��[8�*91�R�\�Q�	��jH�-E� Z�_������������0�ЫI���~�����$m<���u�Mt�VNΰ�ֵ8=�u�S�8���^��rC���چ��ZOͼ�!T��?�KXD�l�	;R34E,d�A�RV��#�=���q	O�J����QY�5�����O�k8�m��C[�>���t��N]*����n�o&��	�P�H� x�6Bf7�4��1b�>�S��>��śL�5Kx��p�?B������:͟A��}�vS�D�BD!Ђ�/*��ɀ������47L��5�VQ��˪�H��gp)�NO#V�O�2��˅L�ܐX��|����S�v�*C��D''s�E5��Ì^J���=�қ�_���X���+l��(N�ړ�g��I\���Na�o��#i��K��Q�ݝ�Zx�x�ҚY�y_���\󖘿g
V�]m�pm�P�'wb�.��M�hD���������#�t�'-�6h:c���/P���Q�DA~,�҆�ք�[6z�>���&}y��`S�� K=�[�� �n3�d�ݎ\3\�q)��z^yvݞ��/vt����ȹ=�����mf�j��i�#��J䁏��|���F[�z��?0���(tz\
�Ne���^]�x"�f���Dkq�M*u<����#wb�H���~Ddcmϼ�tc=�O����RM���A��{
��<�Ϣ�P*}��O�R�6��Z�ĖQ�~���T��.ʩ�^�%��*�/��O���~Q�(w=�p���Pv%4J��(*����W7�K����'Qc�8�n��% �h�φ��� I�ټ�G ����P����
�K��b8��o9p����T�C��xdT��:�k�ſ�(�ؤ%sf6���MUܩ�Cy����}��:ꥭ�D���pP���_,K�fIFW��g�D&�����!V��N�L@:�1N��4�=s8��l��*�1��0�u����9���eD�f��]�J���n_��ؐ�?�+PՉp�>i&���<��#����#-χy�=C���T�
��f�H�(����Xk��)h��Q��p[��шE\|�#���S���'������_H���Z��C��3��	X��:����ׇ�]�H��Q?,c�Ǒ�;"z���u9�~!Ya��3��N��n�z�54v6��h��6�r�F�$��Rr{)�7Z(J���hMr|k��~A˟���i�ڧ�/�%d��t��>�S'��J*�hyD�/}�!>qEo���Ѣ��������W��4P�Oޒ�D�'W�P�v�l�U���v,_�yj�5*˱�X��
�:N0��b~�I�|��%Sz�%;���(�?�[
�����FѤ�;>�m�����)W�0�ނ4�\O\��Wo�V��=�Kl�+ź�4����ߌ���;҆(������;2�F	ɰ��\¯�-��,���t9������AX��H�[�(�]���+��1V������#xL��m�N�n$Sw���� x��؉ݻ����r����@�*�sl.��G~~�_ph��\rLz��i8�@e�a��#C�~X����&D����vdؐ=�?d�3��o�I�s�)GS������_Zο����!���Ap������1H��TX�ᨠ&Z	�܊h �½�)�2�Y��w��y�{,1�S+d����%�\̐�7�)���������β���z�܇ �Yo
bc�v���:	p����,�\W�+�GI��7�O�!�	��R�&��1C�4��|D��>a�sP��Y��">r7AMc�_B�I���	+8�J%�!ωE�,"#�R�~2S2ɛ�=�1��Q]�xZ�~��_b�D��Ǭ3܄��I�$h�l7ޑ�ȯ�Y�08?4,h@�����Ŀ��hm�e$F���ލ�o�H�!K@kA����́���W�v9k�o����Ȗ�P�WD�=Sx]�¸�Uc'���u��Bcǡ���곴��ɝ����c�2gTR�Д>��:�*ܿL��߾F�Qc��ڊn
v�����Ko���fU��P��#Q',��������B�=���Ѣ��_�2���>T/{�e5�ykz臧E;�^�,~z�@lE�����V��a���b5����	�'�������P�t����DV�#i� �D`a!p�[�3�Z��st��Q���ݭ[0U}���*�(�n۽ʶۿ�s��`|���G��������eQPq5P���j
G�Lav�0up8��2wQ"b��&��=�u�ߴS�; �=��lI�ª����uq�1�v�:���j��	���RR���@�tI2ԡk��H�hV��[r�e�k���aE��E#=6-9�=cZ:�� �N��ܓrS�?���F��!��Z�nV�8��Z�����p�����CX[���*SSXۚ�t诤'��<�!�d>���15]$M�vՌ6��q9&�h��VH�ǃeP��c��	zv��x��f�;���5��j�f�
��S���g���m�"2-]��)��4_͖���}���@�(@H�zd���Xtex��l1�3��eI7�7�c��[��"��B��5 [�	�S�@/]���S�P˹�p&6�5
��BDc_tQ.lt0�E������g���fFٜ��L�@�ӛ8�����D����q�����_kDA�@	AE��h�����Q^�
zn�N{����M�zH_��:�F�[���p0�5]#��(&�!#Z�O��~j�V�2�z��/�T�6������h�&���Xy����G�Ʃb�����"߻�U|�ǆ\$ ?	�T䤄j�3C��-+Hzn.=���8�,��8%�w���*�_�ij3Y��Ls�R����<�L�+����y
P��7�R_8Ś��g�o��1���.$�;���[|���_B
���Ԉ�Cጊ����b�熭͙d��2�+2�1؟�Y����F?r��45m���g����gƦr�ˣ���H9�%QCO�a����=_Ƞ�`eu����%�O�vGT�RVe�M�(��N�8��R2�]+�;�yap�	z-��
a��:�O�����]�ࣣ��cm�T[~�ɴl��Ƌ�$�ܒ��P�C�h�,c�$l1�R�]5K��4ʼ�t'쬻�x��y/G��X��� I�>��~E�ie�����NR�Ɔ� D4Ai�i�y3SS��r�-�+P�[K�6�+��SrM0Q��F��qQ%dĊ�RRv���y/_���xw�n�'�WE���^����Td�M��a�$��Q�2��ګ��97�	V������l��6���M�$������S�*���R�(��=:v�ﵒ�u�Ax���]�/��9%F��'k0�r����ԝEw����NV5��R�^<,B��~5��E�<�:B�2D��s��:�1<T���Z�,��:����ϐ,oC�ф��՘;ʨ����͡De3�~�����Z�K� n�Z_�o�ȱ�P�>��Y�vc��Nnr5t�HpT[a�^�|�T������y`l5v����ǬĐ7��1"l�'\Ό>�, ���RB4��j���H��.��7�n޵d7�	���P�{�{q9t��=0d��0�%�A<̊N���|)zx�p���y%����?��r`�ҹ�x��-�z.g�󁈧]��z�*İ:�b
7V����l&;���L�F�v���?�n*��X�m�E O0�f���#D̡K��ɟ6j90�N���R�<�l���n/�|�c�������`���3~`�b�eYv�F}�V���޶d��%�Z�P�U�Z/.�8�*d�Uj,����}⍱��!���7H�oZq�|�8�V^X\&O��Q�Q��Ë��Tw�BF����P&����i+T���c�ǅ�xv_��<���4)(B��E�;/k'��?�# h����Y�ďd�>���&�}�N$_Ѐ�>'m��iAi"�� �E����݂��y�J;�w<;��9+���Z@I�6Z���n�s�i�tUK���Ѩ������_:ڽ�$אd�2�JK~T�@c���	��Һ�|t l�DXL߻M>�_X<�`��ap}��޲�{�1Q&��4�Ȩh�E��������<\a8y�/�mwÃO��}u�+c��Cv4�;->�H;C�o��e�_�	f�^����_21J��(�s��-f?|�m�� N�S��A��,��REi����O7�?w�ݣ�Y��@\�S� �!Δ>i�D��W0���x�<���]�>.��6V*���1/n�3O_��3"ǐ@�H� ���#��5˩�w
SCj�v��l"qb�V��5D��Gwo�^K����LZ�}�g�i�����Ãê�Ei�١2R#�D��oW�/8o͢��f��~.B�9 ��e嘬k]%��T�����K0�(��h��_�6qgY�1��d&˜-�a�]����3�(�~��3�%�(q<��i������1?/���x��{
��u��tЬ��gY��X���8�����י9�ɢ]�/�E���!�X�6��JQb�A8N�h�ۄ`���(*��C�ضs�#�����A'����Z`��<J��cQ|���qO�����X!6��l����ɺ^���}��;jh׃��X)��w���m5�ۨ�8���Ȋ�C�ț��ϵ�Q�e�٢�n���|ƍ�w�Q(�����SN��'��M�2�����m~������O�����5�,׵>��
-ɋCh{!���~��>1ǐ`��1񾩰�N�z������+?\W�ILL���:z��jW�Òx�����
J#���썿��2c��3�s���m� �&��'@�9Y����`k���zmF\S�^k�`��H����V3�%��O���I�Y����:n�6/�q_>|9!��1�PY�_�Y�C(m~4ڵ�]�%�U�YE�{Aҗ�{+s#�R,ބc��j��dU1�����l�h���Yt:�j�Gc�����%\d0�SY����g��ot5ZU*q�ԮO	6���Z�yށg�3���(�$�{B��n�}��?��N�C�YL