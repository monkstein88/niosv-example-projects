��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2i�>�|���B��,<��\ ��W�~��O�?��K��<$џ_�!�ʙ�E�>7VݩGX�& �0����r����Ϟ|�7��.DpJ?
6`��kX+�p[B��,�8��T�?U�� )?�ަ��uS��؈_"�2��4�$�)n��5��JN������Kf������ɯ	�(r�	��sF�"���6�lٝ'���抛�F�Aw��K�C�H�:�={�/h��Ή������Y��7�޹��W1s�Fr<۷���x8OO�٭~� &�����˂n�*{\9�dw��DV�� ��<�0 �r*"L�}E�w=����Ũ���V3_r����x�qD ��E�G��H� ��h����Jazl���m�Ě�_�*ܯm�(�Q9�C�y��v$s 1$fG��a�,�8_]�o��--�	�i��9����4Ŝc���ۃI3����Mk=6x&�>��x�ӂ���rq�$Q��&Nv��'9yH/�eE��s���#0/�v�q���z�����|/���@��>)$��{w�TZ�l��[��Z���t��Pؽ棯�S�P��.u���V6�T���ʖ�h!�M:$�g�Ȇ�����=�yr�s��q<(�PR�q���GF�d��#��4vC�/��
ulZ"����K����n� x&('���7\�%͘�#8�Sa��U�'Q��zx$/�����r���n����*�������r���p˙����X�����S��S�
�ʱ���s��=��s5eG�F���T������B/e)["�R��tR����]�-׾���f�4y��߰d���}�C�j	��P�$��?�6p�1�6n�A|��|CrZ��I�o�p͒�`C~�YR�����t�3W��,��Gm��.�M^�Ҟ��Z�����2އ|�}`�}S��X9�z��.o�L/z�Ke�7(�-����5�Y4��R������S}+ْ�y��^ތ��O���7��z�oO^��_�y�#��v�!���#�D�"�8��ܜ�|(���]��"g�f����)E�R���7>KDL�rh��+�ե�+
f�J��&�~�V�9wh�s㍎,Oڋ9�A����?|uH�U���J��XL�Qn�p,�����+EǊ�Gf�X�ґ��n�s�n^��tvB�Eg���#�����Ė{͚��ap{�mb�ܬ�[�hg'��6�Q�ʄ4�p�imsb\v��}�rz��Bz�Hғ�⼖���a�ߍcf`�u�{�z�}��VA�<K+�z���{���w�p�D׽�K���
��5�
U�mzq.��'�a_ i���`SP���(��#��p^}�P�O������a�t���d�m��T).B��C;.��ae@x@s���9��x�ς��>}r]��;��Ԫ�&�?7-T�6��_��b�}Y�T)D�QJ/Q 7��h�;Z��сr���_���S�������3�,6����Lr���>�cy.ٓ�R��*�L	�?Q�O�A-_�q��7|��F��!o4��7��1�0�3b�dG��U�3fLY�b��5%N���֍�<2ȟ-��ʨ2�S���B�$����unp�3�8��O�yJ����]//��͋���C(
�ȹb���īk��(򂵮�\��R��o�a�萣O��O�������s�����tK-π�B�׫��"6-BI��r�˴��LJ�[q/�cl|��H���>�:/+F��P�B7,p��W,8��8٤��s�C�u��Jz5��l�w���
� B8���v�LVJal���%}��W���v橘ď�Y��=M�=0�! ���VP.L4�,����B��Y�Хڊ/�<+朢��j�Ȍ3�ɑ�/	M޵A�+��r�t��w�����l	�������4�eg�{�7��ű[2�7%cι}�|d^���%CX���֕X�_̛y6����,���B?ֹ���?�u��4�y��ω�Q[cY�H�)=p>�,!�jszs�<%ר$�a�DCp���ר�4�(6 9���}2��8"�&���Q�Y��ϼ�؆@��A2��,W��q��P1!MS�� �$��}L,jT��z�4v��cwe���	�&)n��1j��b��#&��
�>���+�a�/��j~} �!���4��4 ��2~'�2���\sg��w�P��6|��,ʑ[Yf3�3��ְnE$
,~�'�uB=�A�bV�Zf����|�l�R� 'y��,��*k���>ǫ$r�3�<�_�(�?�<a^��x,oS�_�/L�u�H�JB��#�(Q�;�"�-lb2�l��K�|�DiL́���IF��"�(s�}��k7�ց�V��P|�����l+#�IJbF]��d-�s�����ˁ��w�O�$	DM ���4��9�����