// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
pti5B89qQom/PjcrfUj+QraudKvrRFXB9kexI8GCzLw1YhzuDue1c8dwzpBy4eJTT4yvn9RyaaMd
TFJ6C9Xhj9sY6zo7SEi/++9HqFg0LwzV8cm8IAXg2LP2ceLhtqy6Y5Hqw3+4BylV8OV8T0r/Dsln
iFYjiI80bzpciue5zD1U7XLe1goTNNZ9Vj3d49s+gyoyKct27V72MouYIcqjXU4TBW35wPMb7Rpr
d38Vcku2uzLJV0acULmgZrJYS7WxNeiHANiW2MFAMVn6F48YTgsrUVQmH9DhNChZiA5xSFHkcT0t
HuI8IdFRGBTRm7cxXDxqXacc5a8Dk1ZOM5iSDg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4032)
r+bBGpBY3hi4ClXq4a1hWz0BYhr8ka3yOacggboN5YukSx/tlh5DgK6eQ+2Xnfb+V+jNpzRfxyJW
lesTKsADTKRx43oobzZGksX7NmLBDnt2tRfGy/6agQzbGwlolmgLV/OqtISW5BC7KFUxR6zpp9ho
Q9YmT9JddSQ7sucMDP6zmTmSZ5tynharZu19w2WxGt2SqrWgJyq0Rk2cbAXER8MTBWpFUKwJ41hG
NqE9y8J/xM5+bEw6RhWuze3QTM/uxyWjuvLqYe/7J5je6hlbLjyHyT16NP9WRnwct7ASXCCY3WRC
V6WAiaMCXSp+MMZrltQwAWKPG04niJxKRbmpwbWsRlxH4O9O5qkUeX5xJgP6wVJmqZaXJD+cWqPx
zPguMUYG8fvHG/OVGkIlUfOulYf71XcPgcq4VChLrm9sIvUC+5JxEXZaXG20FuGtF8WgOS6Uu+3I
Z5gBRsnywJkJVWy8hMwl2xwG42ZS4rO35NFjwrrgNpHfxSwQ+PLwa5LiUUKb/IBqXfACYqESZAaH
JEpNVP/dJdUZO57MmDpm19FGha4scsrEna0sycOSG5O1Fs1H1YTHVW3gxg551Gi0alSzzY+/lhGW
vn6+FsCvJQTKGl2hb1NtptBljQRt89pc+jL0Fix0CUI9XRsCsN3l9YluRFdLgH7oqRd02WaFEl1/
G9B62j8SuHapoAfXOKtSq59l3sdlhWnibH9/eTRgh0BGDE3hc3p2/Gqk5pH4XWFehSuncC0H+vD+
iUOeVhrdpHPPijs7qHEC7+pt1uKbs48lxoF/3poNBwF35iWSuvMly2WTsH0jqZr8E3UyZsyM74pB
B/wVFp4UVcB+bjnIv48N08+EbrcMsOzcrtq6Qdd8DvjQzZ/XXMi0KwkahzfWVVTYouSZpZ2XFiNl
Y/bSyHIVZa6sHnDKhxgnc04Zi/9GdTH+zPwqKXpnCtLCFcoBt0UDSvezTWVTm36BD0Rp5ebymKTv
WwBl1vujPfm9sQFFAES7EyoXnSZo8cPpqpqMPK1lve+zwLEWAtQYgeet7t+wvEpq1s70rpFof+ly
NwTnc6vx4Ln9klvtNMCutolR1bKX4SArGtAVp9zJh5XIRmqraTd2pjXRIt2y6L4oNP/0rKwdF8pz
5GsCqrHrHzqu7M5chGEY1PO4l/8/HWGYo/Qx5OpdJpRf/qGVGEfAZ+9GiBPSOsOztHqGYWmzYj0i
mWFpUKmJp3spuri7485aFdDqg6QQT1T45OzFdFvh9uBNNWetlmB4iTCPUVk024iM/pCxhS0L92uK
50FR5IiTXTtcvUtHwp51nzDkOfR4E/gqpfdXEcNQ8uF5VKXS2FRxKQx5rxNJRnQhCZo4bZtkRRYa
55LnJ93tgA9jPGGVzRbVE9YaWM/M5Ei5PU9QIZ/m058wQ9fQNtmDgkbQ5nVAfaItJe/0YP7+GIKX
YG5aMFon0GRKdcDvRflawEG3xfViVrhx75pATO/uqxQxKmnyo3BAh+IatCPi4MMEMsKGbQeVPmnt
fC49tLf7IYqdB+LAoB1c2+7Zh+1jHVohTz+RuMZErKo/iBI32j3KlXUMFuSfP3TSzmkhpMxFAl23
PHnX0szMJ7WMBjza9mNmgsYOn/l1aPWQXndurQMWBgfvKbHXA34GPhyQJGovM6Usowlsb7m1KGfH
FwfTUWH0zNtZr9DfJXYVq8Kk+vG23BzDDxzrE7DX2eR0p7leAVa2o2eq4+8YttkjTwIBibKzQDfa
3qY+k22Dt6ZQ/BjvnR48k1HPYnugn9pzK08R7n9hEFGRjim1atMj4fk7rKjoO9eV0Nq+eL584Zq4
01fi/aB8FP4zx0kUl0TIRbHO2XSCweKamiCwoHQarLFqnW9J1Nrq0p9Fp3P7BtLyod1fZBMmjmp2
k4ZkaPYCNZI5TDWDDFoWxR+MXYiaWC+mumUcWQQHnZz+aGR95GNNmpkWlAi+l727ZEcamO87eOzZ
IJs8XDqN+NZP2mKJlpwo5TImvvKj5RACAMJH2poYG3cPa0ThYaT8Sx5zZWPKYnq/fP4335Anekvx
4kveFao3/O8lCswxqLFhObPWxNzPzuAbB+XsIQXVa7tWtcyXO2000kN0ckVmhFSwMsHGl7Uj/Im0
M1/03c38SntKxPIqGaENj8c+vjY4By1B17zmSukaD2uCSZI34nBz8kody7UeiyR37WrP7DOGN4mR
pk3rYK9THf8IZZS9BWV8+cG+NTrUWPSjNL/colaTBJ8Pf5EqEUaIqsRtRb5cRF1+ElHwcO/sYPzF
H5pPQcukblY1/Cvhism+icgzPvHi07ITZ7ZyNumTAiqjxjHjhidl1/tqw+daNce/a9h9VLxxL8St
aV3puIo7+xASte6ZzG9j+fxyzRsxZF8cYZlwuG3GEIlCViY1C8OM+AQHSHNPjU+JPcn8HZuqomuD
5FulTLUje0q3mFkYOVjmChUILaBnKjvKf4a3YtT/AehJblc/gDbwoUIhx6FU0hGOurf7MDMQ0Tfa
AvndjRrCbrtITo7QU7BhRuv3dZIbiYgN1f3iIUbJS2CnySiTDNh4MlkVs6buvr8Bm9ycpCoXYYBR
d+Is5IoD4UDLma/p7AJXdfCTuGaHOsd94jB4aBVAcHFbevL0LmchXtSJx5VV5k+0L2OoYgbXbcqr
ycRaZx6HvnpHfDsm54ac9aaX4XN5+er1zRDQwSal9W/h0fuiWP4+AUxvAxVpBkRYxAxbhEGFA7Vl
0b+bRCyFki1M7IxY1Q1GXIARNqSTKkKtb5LOGKM3z2tLk6YyB2B83EvuwAgusfXSufZbOVsozZCF
DT+sUAjoVfCvWUh60OtZzhsfA3QuLhEOmCsWh+E+BG6aDLDBT9SR4giCkL1zpggSFfL3wlWg30K5
hvMspKUzbo42mUwbvlDKiIcghR8iG6DF+4Piex+LZU+GGFFTQSABFwV3hvIjXswhjF+TpI5Eaw3r
7vpdkJgowiC8OwiLCekLsJ8EgW8fnaeZz8E+/4iY+FJP8fVre2yaPLVjFgt+X9WXkTqh4sirE19y
J2+tjwMdq+C0ICKCDG2KpAUYqvn9NbZJpKcZKuFe/X/F6RsfwfrLJeViB9OORPumcUHgLlaH0uQ/
KJB8uBhXIOyRXX7PiG3KF//LMENFXKt2rQ7YdCGa9PZ53TrM5gdD9/BZv3WqUmPtn8Om9a7G0le8
TVpe3o4tkIkYUc4xL5DFz07xmQ77HWBDWAu1O5+RbRSEp2l3akyKBwTRfyw6LtdDAmq/dLMYzgWb
5esVDJOgqrc0GADhSUz0AOK0eRWFU6Xb/HHF5J9/Hh8AbvauqtKsw/BoDdmem884cmn0HtXnTrhr
pXwww2TJzdnaDnXeK5RglS/+b50+TP00eYCpozWxSTgrKG/M428NUrl0pQCpKgnm1MoEMkCpf4Q1
LP+hfF7XIE2cWWBdEAXE0Oc3dwdmwWDT+p/UNZ02fBE4g+klvlBQbjbbHPsikdxlYORhxZwcWWrc
hz+ExsZFB0aZWxxNi6EaIYJiC4SftmAl7k6aRG+DD0rPKtIlacw7lSOhZoWqiEXwSMIXLHT5Owjt
IWouP7BdxZJb7fmOdNxGSoMyjQwYkWmiEsMSXBVuDaGrYw7+MR4hprrt7f9xYB+UoJhg4WfE958e
q+930qUZtzfwDdoQxqmU5j2NZWMkCNKWlrzaXOzvwpIa+oJrIcNhfu+B1L8cYQ2DM6esmHarkGVV
L7NezXaqqDthjOFB2cKEf1aJCjGlfsRJHMCwvASuJJjOs0LlaIl3kqH8fur7q5zSJ6XHrzLLsS1u
ygj/groPXBOHscc0ZGDiVzvowioDtanuIiUIpHMrp1P8bQ8ZdzPUh/MNhfZy3eQLCYD+pGJqna+7
zGyPnozPm4PI7AbZ65TVdlJomp8jH40BOUZqSUrkacfI3gJYun6XO9ROaJZBrul3lrNCrB+BXIia
WMRlO22dBTjaLd1f46juXJs4OG5+f5Hyx1D8ouUTIqzpQ5GylhGTgGaLf/vmkZgnpLvyoVU+x6yN
otSi0Qi8ZcNxC1avL81Ls0CQeZ4SVMjak1jJAApjG33tr+u0WGlhHqHW3Fz0JOnAiuNkTFUOYwnO
BQS0H3L4yZZa1NL/wI6JaOi135Vgis4dZQ1oXplk6LKhOoQzjik9AGdlBgLDHUwRtYEJQp2kfR1g
phGogZr1PycAqc+AHnGFCU5XSXddZafpXyJQQNhOsl6dWqvVyTJACB2JjbBHibZssCeQukePbll7
FRu6Jv469nRcB8Nq241yUxZzjPd3VIbL3/JPYmrHR6l5dptq4zKjSCzpQ0m3xYSImbFqnrqspWXc
Do4OM/yq4UQGDNCHjVlbQjMeiO017c/VnTPkL16WXs9oQv6EBnOj08iDd3fAUQ4sAFWMlL59oU98
AmYhGibMYKm85u8tLN8tfMgvVJGMc28pCW6POfF+eFK8rT+Wqe/K1c3FDHYb16fIhLSPPCOUjIw/
QZZS3Kn4nk+WMOZ0J7FathtQgI8Xjn1yCzx36G8P8tlxEzMZX6PUTaSTHhk46q48Rf0ioDJyY5aZ
ngiFIoLo2161Yyclg3ubffvJ5AcTG01FdRidWQlp6Zq2bJGt/dgQJQRyMiOhZqrJYHKFrc7Av2M3
AAoduftd6p881LSXaP/Bw9aePGqmmi3Yp7qTxyWJJ1d4Wq8or2PGbR+jRoTSLm0Gydd6TJSh7WKA
aMgwAPNvTn5buld5ic4Iy11UCQ3SXv159e0v79srgugdgxtJN58Qsxtd0MuYPDAdDXziDcYPyyg1
HOWEAjrALepkpXZ22HifDm30N7SOchyNfnB9r8dztEz011zPuzFn8wsGy9DmUfIuFSkSHx4YR4nD
wpa4W+lcSsAUQG17fzlr0fikjsTyIWc29NBcP8fgqsW+akMDR1MoOb7WyKZ8J0L7NwqC2eD7MYXJ
L1jyazQ7Vtdd94dbu9VZvsb5Xb9GrRlxYYNl+fbFKLrjnWndW3dJgozoMXc4iZI0DAMwuNLj0UgV
tc3fskB4Mc+M8slRpBwLtWS5oKiYCN70wqFOy1Mb3ogn1mTd0dNC7FXL1N4WEn7lkr09jCpTM0qh
RRuciaDm0ZM2yqHoEfz08/LxoubQE/8Z6C/JKTbBYIhREzqjKuMr3k761mAiX47AOOfGTYslBOb3
ekMOsiC4QDBoyc9tRI3gLm2T+hcR8k4egf9DlOBXIaF2RdNnEYmHoHueiKmSzilNB2Qc9Zs7u0s7
TAVW3nKQaSB3Eydg940wwyGkgESSrleguemoe4SPYW7rRI0/LoLCF8fX63z+Sw89aSEx+xQSYFU+
j4X3lIjl0VhL1gRhnKm1koVTifqN9UdsKKvp8TZDOJUhJTHmNFwnSouS
`pragma protect end_protected
