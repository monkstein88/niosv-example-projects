��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���~�`���sB�G����fත����y}�e'y5��W�]4>��S���c���,^����ь�Q^R�k�g_6��B��7�jp|&��Ku��V$��8N����x�ܴ�7��a~���0��������?74�&�S�ӏA�����a��!��T�0�&.�~�ܽ�]<[����c���3��`f��"M_0m�_�i2H��4�2�Ɲ��%�qrRР�3�nd�����[���+ۺ�4O(P8t�=E�?��d���NT�R�X��9�A8_τNp���ڏn���a�H>s"=c��8g��8Z��:��B̼���Ƅl^ǋ��m�E�����y�Pv�c݂[���+��I�~Ǭ��#ͣ5+�&C���bNMG�,{�{u��h�����|o�B̌�_���o� J�dM�T��Sq˯�����@,&��������(7D�q���v5qܺA���4���N�y�|h�/�$�p�S~���֏k!�^P)�;�d�!w�������H�� �����KRY��I�c���e�` ����*������d37����E� ��T��f�r1�su#`�Y��P]�
=ƥ)�bp��n�Sc���P]��5��V���>�^�I����<~��BS�	8?���qσ�?=LY�klw4`5>����y~}#��@+H�"����i����a�a82��ʈ�{;�*��S��d{9��2,e�lN��]�S����4l8+�E���d�Ѧ��uW�*�F�L���{k�l���;�
ؔpϋ'��¡��癄cxD�"ze呀�Ι�^�X����-ԟZ��N.e�$���T�X��u�z޴��D�k�u��ٶ���(�����w\q�i���ى�vK>l̩J����<_ώ8��,p;��WSb�d7SM���=1"��l��\��&t�`3��@o1��S�tC#�M
[�I��`��3<6��˒�ʸ���Z\�@�!fgb��-�`��4�%׸�p�Y��J��-�qvFv�� ���G)����	`l7��66I?Dx$�q)�s��o�N�Z��r���:��-uA9km�?f'R����S|��<;���hZ�7O-L��YN�ރJA�t�	Ս���;ZzÓQ6M�E�ّR�pLB-<�:ne�,<�Ih��k~(8`;w��݅ҥ�}q�k���>�M��K�5N��oYW�anj����X��y��췝1=������~G�,���2�3<�=TJ�*�!�,T0�i;+�j���a�n/��o��	Y�Gh�)"2�i�7�g��=S�ɑi�t���|��e�I�Z��7JQ��g�jZ�n�b#_��l$��� 2��Y�<8�����KLUBN8���Td|=CV�Q�����P!���n1G;������O��7S��k@����D�{P[ldli]�CQ����TT���oc<�kO���Ww;�fX[�/&�b�Җ�:$ֹ�JE\u�.{΄K�D'{�;Ve��K����/��,=f?÷�wb3���F� :����6��SGR%�*��v��9��E���@�K E�#[��F�'���n�''�(r��@;���Ըغ��WIM��6��j���ח�\QZ��.J��1Qa}M',2�aIO��ʴ� �c�<�C9�l�N�D�����>Tv���� �9%8Υ����d
�YX[��� xB���v�R
��=�$}�*x��P�<��<���E��Zu��X��N!PkH�*�o��u1����X�n��p,.�ڂ�H�c��Q��wOh��*�3%IV,��ΜV	<?E�]�@�{�Y
����e��ɐ��*դ��+Zr��u��Nj����ĳ�3��{׃�-�"j�tf?bG��~ S_�ݦ�
r̼j��h��a6�a���g��hV�Q5On�@�|�d���͹������ewcIKo��#`�cWF�~ڼ��q�s����K���W�C0���$��s�C1*-"5��*F������4 �$c����Y&uo,��)©[7N�>Ϧ<J&cX/����H���a�������E�Jz���&�0NC���{^ėc����@�D$����ZF�m���.��-f���Ǻz���`���{Q<0��r���%��o�v��b |�dM.�<�4p��ԫt��z��i��4�����5�O��X$Ϧn��.#����Xwش�]��E:�/�<b�+���}5Z7%G����wf�~o�9��f�$勉�l<�3S�/�bI܀�����hd4�����A��j�����F엘l�S%�����E8�M�X:����~D�:0lM?v5/)�4-|\��R[�\!�Ѵ���:�p�n6YQ�?������%5C6i��FUV���Mʾ���U���,��y˅*/,�N�G�l�	��	�?�l�|�W�K���V��a��X)@�o�:�J�M%�v4j]\F�E�$��L�YSN7�]���nT�a�4.�����e�yc��3$݀�G�W4��6`8L�>�z������dw�~��@����G�	lx�>cI���k�<��{���Ru��WtY���fs��}�VN��ry~�4 pC&�n�wY��
O� �S-�����W��<L	�QX"]���y���;�K���ٿ�6<��*�V�ky�
�q�l\��خ��F�c���c�����WnMsU���9���C9����'�Hu^��<�|�~��5��E���"0��?�����������߯tZ"/���z�5sg�R�f�-��j�Vu�
��V��~ギ��b!�30qZ]���w���w�ڨ�����NP`���� ��R6�pݯr����_�EL0�%�y&�ܔ�ؔ@g��UH8 ngsg̩:q��gk�\X��)8�i�xV�i��M������jO�$��@���(��3l��m/c����Z�Grh>���p�y]��ߞB,�?}���]���H�8ݽ�[N?Fǯ9���{���n�B�M�7�*�'m����ϵ`uZ����� /��$�앱��R��%Rn,m,b�L�yV�-�K)��
�lgZ?"��C9A�LTL1S�̈́d#0��k�9�X0!��ߎ.�!HWOڀm�*5��鈇��թ:� W��~��3�&\�$�f	eg�&ԁo��~I�P�e��S�u���&
<te�-Z�p�+4`&��Іhř��	֊���r��m\�O�v�+J2��(�Jz{�B�Vk��ꚸ��:�e��T&���Bǣ��/������w��,HKH!��j�
(>��.�>�k�������M���y�G`d�����T�f���8�
�&L�n��ń���<.S/
�싼Ȝ��~`m�4{�*+鹖�-��0)��d)� 1Zx���ލ�\��~�%3%7Ks
�?��]�8��<,�j����t�����П8rQS��ظ�!��|*܊213V�X����!W��~����z��]{���5k�]��;��Y�	mO��~B��F�1�Np`�Z��V?��]h��o���ggj����9�m1��$��7�m�.�Ǌ:�2{�/lp�׏�4&P��Z hť�7B 0	Y�3%�Җ�U#-< �r�>��yzd����������
��C��_ɼZ�i� �N"�S����y���j>�@����	���S$�=�&3[?�t�T�\�l��[܊+Y�d����3y���4up���VK��7v �݌1��}�;w׊{�Ǐ�t	N�׆�ȶ��"4����&�<r<�p~�f��b/p�9 L�-!�%Y���P��1��78����R	_���_l�j/��<y�V��dŌ�8�}�@-qa��@�_����Ҩ{�����j�h�6Z��@��C���Nk\͡���1	��JU�h�&\��FW�}e���O���놹A���7��C��qy�+��~v�1'�{�ޘRG��E,Os�� �.G�ܴ� 6L����jP�'�<4�n�^��#���C�*Q+hj8������!+��\%I�:�4o�OL���R?b*����n9#�@t�G����9*I����م����@�[�_@ې�꾭C�r#Mߵ��
2�l��ϖ��d� ����M��>��z�!�Y���HK�G����տ.���P�������3����$�\��:	�CI������gLU`*��o��o��7p�̅w��� u� .˶�z'W&M�gY[��j�Nv�|�-�� L��<V2�IfM��e��X	�����,��pM�/�_�j�k��)���������\��kL����9P�k����� �5%:0����G��&���+��CY~*~�e�̶��9��7���̽����Y�$��&����N�?PiY���D�8Nw\#e��T�bx��0������zl��������!�%�L�J�v-����B]Q��U�$�\QńUM3�y�;����%p��
��c�-0��0%�.�+
ΆVܡdxxU�D����q/Kx������"O��qk�x��U�'Zsʇ;E�*���'�tb���߼�%�la0d��`�@<�;J��(#LpU�h9.�,��7�2���6�(Ϫm�D��N���p0<�Ļ�/�����1�mwG5��-� ��us�k�.�7O����bE^2�Ew����V�(h�@���֔S!�y�LRfl����ҦKn-
�9U£�<<�(tHRhcO�W�y�
&�cY�b������5�� �wJ�9�!:��wŹ��T_Y>E5.�@ _���B�o�5�iR=$s ˂na��Tve�+�T�=���=`=t2�t�${��:8B4ܘ�3�7[������|PL)�oɣ���Ȼ:,��**Lޞ���l�c!h�;Sp������nn�ov���%����!�^m�!_Fڿ�je\�M���Mt�N��L>�9�ۚٱ"�ũ�ɘ��vAz�?z���t��LC���kD�;"-%����� @ rvJ �)���Y�`˕r�S�X-��:��㕹,c��Q6�.

�O�S3?�9�7l8���v/��̃>��r�z�8!A}�JƐ+¼G�P+�CQ\�����ˣڡ�EQ�@ݳm$@�樵�{נɷMP3�(R�?�u`�$�KA��Xw���ZZ�h�V`�o�uN��o�F�������fD�X	�#�.�f��Si��o�X���LJs|Cr�]L����$���2�+h�mz)�
?>��p�I���h���C�C|A�?�.|�[&�Ŧpُ@�n�	A+��+�",
�(E��X!��2p��[c��RʓC��Be�l�!���,�Q��H�ԉ*m�g�Rg|^]�Wa��W[F{�g����!5>zD�
ή���[ρ�x�ka3�&��R���U�;?Y����,�$`�0�K��QL/�US?���e��m&f�� ���5H�є ��� ���H�텑('?�*F\�G��	��!
�"��g$Ԭ��Y�a���YoO�������\��E2q����k�$@�A.Ĳ�ץF2���Ȟ�z�������ہ$G��Tr��s:N���uB(�L
��x���Q��vi/���=��(L�Ӏ�x0$t��T��-G�KK�K�0�\_E\��5/��8Xm�ї�<�LT���%%p;��F<����f�\j�^�^�?��,&��Hf�MR[0@6�>�JGm���%��С�Dŕ�EV���	-�WKZ�l���;���4�[�l���ď��h�-3ͳ{#-�f_z�G�'�7q� >�2q/eS��g@&�]x1�P�Rb�����5^�_�WQD���sî3�����
�cV㔤��������ފ�ۭܯ��P#3v����p�o!���t�>��rrH=�.��Hȇ�i4����印��)&d�8����u�;i���5Ͳ�TF��� 9��7�����m�����R�$ŧ��%����7��OBQ����5� �S����a��8�2���R���'�rU��a�;���O0�\��R���#�����`��r�$�r֣����O���:�4�Iym���?o�	n&��������������5�!����ZN���1l��p.��+�E���爸��f�)�,��ie����h=Љ�Qa*����n݆�r�E
�?���s�|s�}�%��Qh���+o�����Y�,b���Bi�X��� Y���5�7�;xd�N�٥HZx��X*EK��)���5m �b�8W��L��%:�d�99�J]"�̔C|R�����y�v�a4x�h�y[�z	�=����}*������.Յ/L:֣�C��¶�e醳�k������eB�����DrJn4�3�Ԭz}�+J@�@-2�>�Ϫ�O�K��ߏ[)MK�	��DQ�%v�R�	D~��/�Fm:D��}F���N��BR;� �t-��uE��pQ籎�=s.���-��x��ˉȥ;���$ǭb�V
�l�Ķ����;�Poh�<�|s0`z����i�n3 �PV��u�V�G��[A���A�9�l�b>����ʞi�ob�ԧ���쪗[M���>Y�q9�{�ך��D5�%�kݼ!����I��Լ=���2\T���L�X�B�-D��9�p�E�hi�dL;8�Ԇ���^���Ѥ�6O���A��^�m0��R"�D���Ϥ�j�=mm�Rf��rG���z�υ!��Q屟Gt��z�!h#���'��}�֪[�M�
zdf��m���zt�jc@�L��G,��Motu�Z��:��"vpX�E Uw�8$�����G����P%��
�8��rkf
9��>�WxDKcpaK{��]&LC��>��a� �E�ܚ}�D r[�����x�HH��/Z�\�)Yt���rb\ݶ�|Q�P�-�`�3&.}�HL��Ӈ-ቺ��k�]:N����"ȴ���
hwO�� -TFwݟ&A�]�8�����g�Z�Z쬾���{Q�8w]��A�Ž����]�ٷOz
Ǫv������NK���5���f�ܬ�➁���29iD��|�_Q��DZ)�+��ݫ�*u�`禗��p2��;>^�[3���{e%I��n�� x;�(�!$��?+v���洏 ������n��0}8�v�m?��K8 uY��=��s*�:M�������$H�o��)G��(אR�ᆲz8��}{� ڊ����?��6��V����U�,!���D�����A��;/\�
{M���{�ba5�th���6�'���b�G�u��߬U4���;�T��fٛ΄{	2�#@�S�f�'��-CM�^�ŎP�Fm"�ۮRY0�y{��e�׵��;$bb���@�*z�U�a��ad� �%��t��8y5�y��Pז~<��ȷ����/;�m�s氮�&��j�N|c7hό���ўF۬�����F�u�(K��'�Gn�1�tQR���1ʻ �ݠ��I�D 1Ƣ�	�fߘ�g�`y��=D�M���k����p׿����
H?ܠ��ʐ�i�q���NCDAM���Um��o!���-.�� X.I��1��5>#z����a�< [��Qo�ϙ{��[*�u}.�?|o�R�Z�\�f{����*�E���Ԝhnt��>H���V*|T�Zq5��"���_�[�Z�]�Â�J��X�{�=��䓶Dd�C|П񊵞_���1�$*pi@v�-O������Z������)�o����;�p=1^�W5�J*䇮��F,}ish@� �Mއ,ַl�4�L���A��^�pG�l�%�<eʔX�p���6��蝔�E?E���V ��:3Gu*���j�d��5m�qȁ
�;��(0���E����&��h���Y�����\~����r���&�FD*�uX"��|�6��T/1(8�E�L��'����G��n*K�+�̭M�Թ��.�X�N�u�=,�~�oL��QsJ ��o�$^��_B�c߱Q�3�V�0�'򙡾"����L�����8�D7.ݣ����ă���l�bF2*��`��T�}{�a*�N
/�鉼'j�6'�iX>���e߽T�h�����[�%fSm����Z�����íe�b,T�vpf	��&�׳���5�p#���OGr��HI'AnD܍���%�.+�Mr�NP�H��.(H%,�?�� wg���$n�v�Ǥ�^�q�{��������"��	�+3.r���ԻTr�E�%����V\1���ة&��Xd;dsJE&a#�@�beY���!�la,_?��v,�.���e�?�xD��(� E�$*(��I����W��J%4PT������GW��V%�LoTD�%ج��/(���/A�Ŋp�rv��i';K&	s׉*��J�M�1Z���f|�U���%�`Z���2!�3�E{�$��h�QꐎDO�F���}[��[\k��l��#D+b��5�n3/Tףo�H�B�����+�'L3ɪ"�mQB�ʫ��f�����yV&��G��h�L����
e�u��[U �D��s0Ji�a�.�T�Og�y-���+Ta��0��RG���,!���+�`�X�E[3��t��I�l�����Q~j���$oE���RĽG��g~t;Y6c��_$Z!!�±��$'�6R+��S�&���3&9X�����4w�*���C �&ʔ'ak�@#�c���a����y�l53��N�r��;�����&��]��4�P�L:&/��f*\�>F6��Sn t�}a:X���6��{�S��l�QK���d�����#~.U�fl��SXIt���vן���6�(��t�
��5�8Ũ],�5W�x�&�'��Ã"��ʪ���8���f��U���|�@z0l�tos%��x��w%���#��0�&��.}�+�ê	Rd����_y�:,��nhm@��-�-�q4�q��C���V�u}�7M�#P>���EI�+�*��%�a�r*J �9��c&K6I�=z�_t.��=<d�8������X�`!b