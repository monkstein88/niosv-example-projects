��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a���V�h�x�����>�`���o��藶���ý�T��U�Sy���So�x����t��6T�0pnn,Y��FJ%
���t4��b@�3|�W�zR5M'�%�+�o\n��m[��v&��N���n3mŅ��}L���"�̞-��r��8tHY���� :�.Z�K���#G�*�5��s�e��gl0I��ddY��ܤ���?�R\(�n�O��6�*y$�����@����1Q�;ǀ�^2�a�Z���G��92΃ 1��+Zq�������N{!���*�)}�te�E��|�N]G*�۷t'M$�C_g����|�yAa�Y���eĥ���n���2�������(
�33�Ty�V�)+#���f%	͸4�Gp����v]% o�� %�/k��O`�����$��:/Mg��t����e�An�U[�D���n��X�|$�y~�͠�����e��V~?]g��%;98Sm88�NK���F��d��t��9���t�Y.^G���HC|��:�B���Շ�f ��Q��!>���O��Gp�n&�i(�ͽA��#mq_Cj��Nz>R_�R���׸q:]� ��VR�7�=ǰ�)�)4^�4%��>7��O���os�Y}������\#t���sS�2�"�
����J'���Hw�}3���:E���ޑ;�S��)�	�7�ʹ(�����}ƄQ�������������Pv%T���ב!�2�����6��`��!�>ӡ,�EΔ����D-)�o�ha+�"h!�f��g��A�k0�t�M)�/6+=肇�YjS�άW:�#��T�{��vp�Z?^^t��E�2#6i5H+]��Vo_w���D�ް�����"�-?+�d�\"���ؾg<�@Y��`�-��Ǩ�񡧄#�OB~{*�o���#�\����Y	��a*�}�	gqa�|b�]�D7�Dμ�V:PBZ� �JB���'c�~��5a�G�<�=�{	V`�ͥ^
�����'�|t�CV��ǵ���a�MY�p��S�f݆����g����I�_�����)%@�$��Z܃�1b��M�6��7z�$c����p�U��I9��������;֬���ؖ�����
�;�'B���J$����Xp ��,$,���Lmt�WxVfv�����AlM6	�p=�%��䒝
��Y
T$f�a�d�qf�p2:JZ�ջn��� ��ƺ�ϳ*nsN�O`/���ؑī;���OQ~��X>�-�'qB���ٜv���֐���D��'�Q���8�c��g(.S�;�|�a	X�����%=���_�iG��UN��O�*�C�% :q��T��v��4�Q�$��)�K�o��5�d�R#5��2����9Iq��;`�����	��(O��������C3���x/n��۳E��-Fd���'���_�H��g^�.��뽗r�ǎ�Cr����<4v�9s�`ؤ�t1�~� ������h�%��j,��l��Fq�AcFG��ö�y~9u3T{w�7��~̹*g��;8��0�[��wMx+�'�p��y��ׂצ�Ku4�g�<��&��M�):>������9�{wH_ό��I-���3nO�ʝb��yO�U_]���w����S��qF���up��h�uh�}V���o��zts����ƙ�2�&G5B��a������iJN���sJvc�EN0H[Zt�Y��Į^מ��ǉ4#T'���Hs{1h%�w�����"���Ó�z ��v��B"���n�,Ȏ?i&DEqTe�뿼����uSq\3fW7���ޛyb��|b��ON
�^��t���Caa��������W7��C�9r�Qϻ��MI���|0W�v��ΐ�����GKV�Υ�ļ{���\[�79M��`�G2�0Púq;4������,6�.Rc��3�7a�R��)}�}�8h�j�#� )�d�V��O�͞W��+$����8i��i-��� c���|_ReAF�r;.��}��IB����������,bϩ;q C �W�O��� ��������ή'z�˲�
�F��i�Q�����c����hV\Y�r�,Tt 9�L�r��X`��E����g<�2��O�&��s���Ԣ�A�*9$o'2�t�ɇ��������c��S��1�;.��kPY��Άd��u[���h�BH�euً �b�{'��~��S���W�I����Wxy�~%�Cy�o-��s"�����62e�����߀JlB��`�c�c���7�਷yVWb��F���О���R���5�s��KT���x���S�C���O5?P�lV�4��%��o�oh�~L�{���~IP�@aBj��e	&V����4� y ҂�9ǘ�9j'c8z3�Y��-@��R�p0ur�rB�(�tF��cLv�C��B� �o���Hx��ή�[��.�+7޳���(;)G��U�@?a��uʊG�+��py����TcB�<G�'������ws(gۚJE���,�y��F�=m(��9B�5���s%32��v��~$jmeV�6�r;$�%E��)�ܴ�D�ȸ���RB���T����ĳ��
�S�[�q����s�	�s7���W%ȳk�6���;�����=��xXh8
�.	d-繆m�wZ^� �s�N��s�$��,*�̥�YU:��g��/.M7���UH�ӏw����\	��xg&bD8�q��L�lF��1P���0�j��:륮,�δ��f���-�!x5O�ei݉�Ʊߏc�I�-,+�ϸ�{���Ũ��t�;�(��#�^
��^oَ�����ӭ�i�q�*b��4��^�q�ݐ¦�]�쥦�{��� �R��F�!1!R�#CNށYIm����8S ?��C�7V/�Y� aS�M��	�ͻ�@Lf�ԉ0󑴳������<=�xV���s��+*�~�Ao@�F|�!v&�zv��bT;v$�J�3맳��y$V<"��k�Q�`��J>	�&���r���S"��� y�����bY7%�����[�[� ������a���Ʊ�fw�V0���c��.�#����F/OS2W�Htϵ���;�-�2F��}$��GzDU�j��?B�S���K^�¬�h�,d���fq"%b',�l?r˙��6��3u��h*U�����\��|س?G9�O�R�d5x���u���'�h6�RGJ�l�a�]�JI����r.�Z> ��ђ�@@B�︽,��<+��I�z��lԳ�)��QD'm�ɀ^g#ɝ�G@R��� �@�f�N)�
'r(7"���洷��~VO���s0�TDu����N@�U��ۦ�"�VG�_/L��l�^8qJ�&?�3�
�J-�ϱ3�z����5/�Ε��`,��"�7���݃����?$�C����4L>�D�Y��t�	ͳ�ʹu�����y�5@M��|�Ԧ��Y�g	h�Mf������Lt�����no(�z�K�fd�3� 1�`�����cQM�������]k"8�L��߿U Ǝ�Ncxw1U�vp@&CA�*��,E�oޖ�;�k�.����r���n���M�^*��F�~�U��}B,�x���4R�toY��4��.�UlSئ�@.d�?<i9�T�B_aN��5r�y����2B�&�;y����m��A�t[�=��6�S�\\̹����zX*��o��L2�X5���X0�l��C�b1�.^��U<9��u#�)i#�������m��K�,2x�y��Z�F�4�[
������!���hJ�*3�Փ�BY�/�ԏ�>�8/�,��ԣՃD´hJ�VZ�Bn��
��.���O�3v�A��5f��a�}�ۈ!i���!�#���N�Lrrb�*�H�܌�%��W/�ʘ��8�]�o�=�.�an�;�[�!PZ˴�)���ߚԶ�߈OƚQ`0齱��z��E������u�ۖk�	X<6�<@�J�)�<^6�3(��v�%V���,�����H�K����"�����������2�B�t��p������w��V��H+��4����B���܁��� ��$�+�V���(#�u�����Tq��n�����+�+���ɺ�����"ڃ嚠�"����`����-l(0���R�ù Tjqf����9����i}�ֳ�]�B8��̎t�"l��'����V۫>��k.낝��N�_
*�� V_����k �eDK^��a5��x��K��zA���M���-ɧx�����߼TQ�+�bs��7t�} �Vđ��Ҕ�ʀؕ�qBU-��&,��k�X".xk�%<����}ҷ��<6@�C��k�䶤�n�?f����H:����"l�9�U]͆��a������T��>^hj�D�؟Y�
�R/����G������t���\%-�K��Z Nj���5�`[R´l����{f{eR��E6�RI�0�z�����a�i�3���d#�R�]�i��[\����P�c�i��m�[�U +4�AZ�� *ޟ�J�(�(�L|PXd�!˹{Hg�v��M�yN��(%�*>!��{A>�a	]�\O��	��c�����.v���V��{�{ׅ)2%(o��˽�Ri.^��wԧN��p�;�o��	�
�]�������~AI�T�:��.��U<n�۳U�d���Gp�YuykG���*{ ՙ���$�X����ј.�^�8,�ĝ��+s�X
��;S�A�>�i�R�+��d��7��)��٥k~QI���IC �ū��3)U�D�i���3Q_�")�ϡJ)���]Uh�0���&����Hl��)��ׇ�ۃ<J��
^�{��;��OV)�s��ɦɑv@G2f���v����De�mZ���Did���@��X]^c�ÁP���S?΀��-�ܮ��:�6�x-!=���1���g&�x|m!��G>�b���Qɚ��u���;'k1��eA��^�$������*o����?AǛ�16�`�/�%R���pܻQ�,H鐑b%�L�ߨD��D]z%R���vo:Z�Q(B�$ZQ��,��.k�''�~t���ƃ�Y6��+��ʶ���םN��&œ�׀����S*�)0�KE�:��X�:��<�p��K�"A�h�Q��

��o����	|��zl���Ȅ��q�vbd{�&R8#yCô��=]��v�`��~}�O���a���H�����8�$H&^�	˙m�G �傱�`�(uT�u*��*_�3[���2��Ï._�n�3(j�ih�浐�����G2R���@W������o���[�h���Ǻd_J-��qY���qn��������$���k�t���������]M�z�R�c��Z��L,��. m�,}�/Q��sJS:aΖ������p�d���i��'���<q�GvO'���b��-��Hkٹ�-�����	�#�ҀaM��6#���i�� �eA�3�H��0G/of_�L�� �!E6��Y�'~�\������+�䗑�8�8ǹg�_���%	9�J���x����ЏIN<��С��!�Rm�T��R��d�϶�~����7�Z�t��L�[|7���.�W��@�Ӵ�g,Ȟ�J]��`졚{��d�]W���@�_A'/f��'X�8�/�{�]QS�?ژ��<���q��{W�d
6h�d��>���@��@H��#��`�(�p�>B:��mV,5�����|-2=�{��(/�vS��ǯ���"��P԰���23��D�E�'�����=e+�(����#���� {Q}MR@9"l3��o�z�|�F2�j�_�y��0�Q0����`������AS�{�g����
��x��k�����B��V�]s�v���;ƈ����;٤󥵡R����~Lcyz�S���.T�)ߌ�32Ѧ��#�:��(��r�=`��ʿI}�#��J�鬵���~jY�h��ME�jr���W�{͘�Tm�m�4zC���>�}~��y�԰���tq`w~A�?ɓ���1ܕ���������ɥb��-?��)�0U7c�����B@�y���6-���@1���~s*��={m���-$�Sg(m"ҥ��}������
���F�� ���c|۶z�G����R�7��������Ƽ����E$|�m�N�80�  *�������!�s�it��؆��J�;̋;t=�3R�{��X���~ďF�|�NL>/2tV��y���R��9�Ҫ�����0���ge������$y�BXL�'�22?Gج]�휰@\�vY�������!�P�J~���_#K�y+������G��qQl=�Ko����Ω�d\��+��?��s��"��ho>��N!h˷��e���Tz�o�G����rx���x�X�̘|#����Z1�܅�)�^V�n� gxx�Yz�|�֤>���]�hDB`�`�j®N�cmud>�S��4�q�?�=�.�!���[G��zA(����`��A|����|���z����Ej��L.�����gWEp�>�XQ&՟]#�I,-�5&�� }F�*F?A�����3�O~/��\	�ȗ/ʢd+�0�|�}��T�s0��U�u;.��y�7����yd�ԥ2���%�&�D����/t��rC���T�w�˚�o�����E&�Z�3�.#K|�Nf��J�:�Nv�E#q�<xY��� �b$�D+��]����ۄ����|��&��1^o�h��f�y��{�tջ�89Q쇑T���0bM����y��&<e36��E  �l�fw�����N��k��-ª)�p%A����ʣlH�k��}=���(�)�7R��F[���(:���mB��F���ߙ`���ד.%�
QO��}H<	--}���\��X�h{��wZ�
2��q��Nm�zѓq��<A0ćkh����Q>n� ��z�q9KOh	~C�a����j��f����h\ (��
���l[�I�بFU�	ދ -b"51�K���9��Hz��\# cD� {�&�@��� ��\$h.;{<�E����5ޟ0��9z��.�G��BB�H�e�E��󘏙�ٱActS9/�M}��2�a��;#����lc|�2���/8����8:�_�O0��ܮ	�-)D���%��Qe���N���?�"(�-l�
�B~<�}Ƅ^�-XTi�A�P��3���kA���H��d2�M�@ͦ�)Z�{��5��.�pfn�'�@O5� m �`;���eGV�"ѣ��CC5�I����O|������"�-��0}Թ��5u���.���P2�Lb�hllb_͓�����n�S�o.���A��apPVA��,W'S���)��p<�?�|�Ȟ���"TKq<ؽ��='&�s�?��2c�2)��zd[���/:;	��7��gH1���]�!@�����l��ЈA?��o�& #�S���AT��u�Th��a�6A����+�_v>Cp�U�B4
 �G�\�X���DR|`�)NQ��=4�p^QdK,2�-x���@���1ي����/�x���]d���hٵ �b�R��o�<Q	���6��G���&a�R$h����\�K��>�q��w �7���GOY1Hw�Ɋ�nʓ%��g$�ma@�k N�s����ʶr�y3<�(�V�3s8��k	��f��˫Lb�s��&XI����ﵠfR1��7T�����2�N�ۦL�JG$���f�x�b�	,�������� ���-)+h:���	�����)��c[b"v�E���
F�P^���l�����%yό�}��h����*
:�nG#�;|�N'��X������Տܼ��O)ђj�2�w���Ѿ**:��=��Tqw�� �4��6eR�s%{2��"ѼU�|��|� g��:�d��/�@`X�oM�w\~>��L��?��SJN��p%Vj3��&X���,��׀�T�o�#�0�A��KZ�et��/'�
��f>zʘ�2T����O�2�,�t|��A]���3Z�����K�����v�M�G��#+��'�
<]"��ŷ��c,N�~qc�#~���e����O� S��4"z��6~���+�#�J��>b��4���m������죢"��9�-`�X�Lu�,��)�A�
����Q{z�{n�8(	Q�Z0 �r�${��L�������#'%���Ɍ���:��	��1��3+� ��EdnoVf�ȷ����:�X����� �P&��vq��f��fwm�|�O��?
z2���<�˜��r"��.J^7�Zl����fuݧ���i<o�P��@�di�!���������t�sҩ�f���#@u��D�|�� ���N�R�6����N�CVL���-�5����KZ�3�S.����{L�~0��X��i�_`��6�i�
��Za��#*"��ƻ\q��VC*G[�V�'�Ey� �1'��3o��a�̝<������'⇚"�W�1�T+���m�CO|��TC���/B;���c��޿w ߩ����o��@�ahQm���α�wK7pѧt�����E!_� �0��)�Zo�'�qk�	����r�w�ˎNJBPtģ��)��]�G��9О�	��,��^�Y�VՓ�@d:$�M��L�IZH ���nJ/�M������r�$���S��D��4�h��/.ֱ�A���ʶYAP�ߑ��Q:��l՛�!Η�z!������m�ǁ�Y���|ɶR��!!�l�-Գ; '50����\�W�p��}ݞ�mA�9(�QP�qT�������Q`�]���eb�X.o-���u��O�-ၱ���r�Ȫ�f@b�6�������ّ���o��d��従�j�N� �Z�!�p�Dq�ڸfd������~�_6f�e��ǁ��tv��3��1��+v6��%=B�@F��E�4;�-�{5������sT8�·��d=���(���`�*Fb����^�� �U��v}��hLa�8~��|/�|��o� 'f�&Z�iʏ��}��i��k��
�Q�^F�ǽy�Q�*���%ŖA�B$F�MHgS.$�X,��#������؂�.? �(���I_�S���̍Ю���	{��s�#b؏�� 5� �t_r(�{+ym���Ag�&@�#�2��i�������BV5�cO��X׼`����4������U,�R/�x?�����ٜ�l�b��6'��ۼBE��//5S��y�c_+�D��hd�eȫ��o�Lρյ�z��\��.ILf�Gڒ�@#�>���ߪ?�
�/��vv��G��_8��ư$�zU���w��I?�<c�D�R�A�kӯZe+f�=y|K����`Ob⼺颂_�w�j߳t�����m�p��+iA@D�_7���~�|�t�S2�B�f�>*\�y���Bf��H&P�S)�	 ���Nb,��|�Ӥuͳo��F7�9M4�f_*l��[����B��+��mrz ��e��ec��CX����M��i%6������<ܕC���؜�}���^Qo�U�9>N^X�N(P�LG��N���HR��`�[�,R
�/V��W�m{7@$����;9s�p����Dp!ϻ$� ?e��;�)	k�����M\��~�� ]�*v
���X�*�x3Xb�O����1��|����q,;�B�������;�D	PO�2[*S���, ��*k	�/��!�AМɰV�H���q�Fn�\B���N��x��qQi�� g��H���:����̄� ����~��xT�PH>,�JH��mg��W�\�W\�I8w��[8�Q�Ҹ]Dϵ�j�(��WƥG�g�X{���Y#x�-�R��z�(Х?8!����^
\�O��P�