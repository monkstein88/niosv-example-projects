��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2i�>�|���B��,<��\ ��W�~��O�?��K��<$џ_�!�ʙ�E��,�?�����2P�i���Te�#S�յ��-�4>��=���c��-��6t<�g>a��{�6��ŉ���%[P�}�O<��d�!̫��]��C_p`&�)JLؠ���Qs��/�Q|0���6U@���y)W�ſ�N��~g�kF�����B��Us�n�Oxӣ\X`�M�9,ܸ0���Q��f�A#�x��f5�n��i�j�==�:8��+�Cv/�2-Bo��JZ �.��ވ��-�@̲V"�>����>Wb�����
^�Cl25�������[sr#���2����+�����{n���H�:��r�fGzc�M�-�j�d�ư�5�΋ˏQ)�
!� ~�p�F��8���̀��x�P
�z��䔾��Jl��{N�ϩd�׺��&�~�������*F�yX��X�q�{!�S��jρay����G��eNE.# �dB��Ձ��ʋ� �w1j����]��'iȠ�|��LZ:ɍ٢,�on��=F��"����cEV�,/��\��6�{��D�t�������
~�����X�|��u�y����F��
�g��ťX�K~��F{õ;�}���B�"(��X��-�B��PSK���![m.| S�1K���yС��pa1p��/:&d�/>N�[��u�N�����f�%�!}kW '������@��v��71�����Ѐ�Y��}?�N%��#��`���z��a���YrZ�
<"�M��n~�X��'����THW�6�}�����w;b����t�N��_�oq�XQ	���mqoH���&��״�ۄ�~���^��C��e���=�����?������r����flFA���~�f>U�~E�2�֑�*v f�3�������u2�8�6�9H�=�9V�>� !E�r���
K=x��R!/b�bX���	/��m���1Y,P��������ij0���F��	۠�i4J���u��� �0�zP���#�T�s�Q�D�����E"�񥇚�4}�B�B�������Ʋ��L*�H�v5����MݻS�!�H�n��J�%�-o�$�����Z���I=<3���Ë���4�ڤ��D?��T�9"�"�e��y|������[V9�:ЯO�I���ܫ���n�F:�'Bش�A��"7���Yc��۞&� 6���[*�QN���:�ԉI��@2#h������{�;���Q��Ë��1��Duy�f�m���LH#b���RS7�V����JV�??�z��&`�Ν�bA�Lºf��ف�87huٴ3��DƦ�f^��Y�������ci$�/�d!�aH6v�:�p#�l:�\�ĭS�y�=*H(�P�<��y�1+9Y�0>U�ڒq���J�0`Яg&۱S�N�vL��~��9K����#�#Wp�_��uMH��j�]��*,WV-��"���\e�%���2�ŌSl�߰$�Kf�J��!�7�!w��-�t�[�����{A.�ߢ�s�y��C(��	4���h����'�b�y��E͋H;���'�v���[_ �I��+��#�S�X���E�02�17f�1vēPV�vhaHpYB�A,v�H(����
�EEO@�q���:���?�!k��e�	N>��ĊnyZ�.�"�6�	n2tR��yV|cc�D�J�G��;��(�Ȗx�s\e�۟��p/�M+b.����[rs �͜�f`3�Qa���#n���HL<�T೜�����K���i�4�3�ќu���Y�Ƒ0Q�������}����yG�į� ዏ���U��������q&��L�����b��-�3Œ�Gf�cX�HZ\o��}4�h맫H܍q��l�cU�>��p��\�G��͏�=�W����C�0�1]�ūY��Υĩ��SR�s����*9p�8=�v��I'�7o�����x{G ���G�7������V�U�WPuK��J�	53�	�����(Lw���.*⻟��J�h�El5_|x��;e�(��**�0Ċ�s� K ��ƹU{�W[t���i�A@
�����f��E&��Ӯ(~�v�F�R�Z5�M�-$��2����Qޏdc����G�yG6P��zl��9%���BYJ��V5"�}��#�߄�C��L祱��'����(�a!�.�T��c�����B�7�B��6Y��d��xJ?�������Ȯ��C���C�b��D ��{hfv��0��W�b�h�\�̰��8���J�t�y)�lk��ٮ�ܪ��W�;��W����0 /~��~�6�pN`�NOux�-�oB�z�(kі/�]݌��?Suo���(mFt�Ą�o�GKAdzv��
aU���u�&J:�~�~��p�~�����a~�U�r���\ �J�n�Qʼ�����.����p��
�,J- �xQm��׀.�+t8�pV�պh�`E�� '/<2�d�rDAr�2��R�7`P}X���d:2�S�	5e�P^i�����{�������(��&�����&��Bb�{o]�;�4�H߉�T�Ye�W��}2��}�t��a��@�J#�fa�w	^�Ԟ��t�IT~�����3����y<�X�NOWeS��i;��T�y��q�߆7`.�4˰fS�e
�}����?9G�.�.'b�Z����g��g$�N���d��{���+w�c����E\�d8Z�.EN�%� I�@�W��M�f��nί�S[P��Y��25(�wI�R�h����Y�wM|r5@�[��:d��� �dE�Y�%90p�߂�h;�B�Y���B;�J;�H֚q����W����rV�)�qt��M9��::��7dڏ|�5pq�\�֐X�F&S��=�`7K��Kca���v,'cPZx��3.��4�!�eE����Y�d�4XI�J��.)IL�)��'���͎c�s�����9�'���\[n�L�֚'�Go����H��ڛC�I�e�g�����P�W��Ԙh�6b�q�`��G>�y�����O���c���-��k���>�(��2-a��iS���C�Xr�^�h
���?��I��V��nDΊd5"u����q)�c@h�c��ɳl��d�2Z;z�0,&8J��?#f�����z#咯���M�Q�|�+aZ�E��U��u�i��Sa0`��0IP"�Fy�u��n���(��O��8L0�i��-���#�����o�9���u�7?P���N}��8d���e�}yp0"Y�YO�m8T�%�e�e�WX7�I��ض���u����.d����]���Fܕ+D��j0��=�%����J�d��N���L���?6��mW�x��ȏEF�}">$%�&��T." k��M؀! �5WGe�gc���V��4A1p̪������@�:��/�>Si:-��-�f����\�`pm�%g�UGY��N�k�O�I���d�|E�21[Cӑ����p6c��j��b�v�O�=W��Q��cA1��_������ӝ�S�6tǬ�cTa�Kt��aֺ�u���h���A��*/���n���\�Il�ٻ`���r�֜^�X��	5�P����=�:�5{\Վ�7��*��s�����#.mS8"Ke��I�3�#��L&w�/@=g��-��_=�)d��(�9[0�^���A_x���JV�/H��D�Ė_�鎖�2��6��'pU?����'�`�&���#���KPG�C3�����\n�Z�P�Q���Y02�!���w�)��\��.O�s��Ԕ}̷9�fH��Y�!�O������/�:%~u���H7��S���p�������`�[�(+���|V ���Ndo�����҃�Sh�n�*݈G����W+�����^�d�cVv����A�]�'4�3\���NI;�9u0��!-�ȭ1��*��Q5O�0����?3���85[`�
J�{O��*z�(kӌ;�Y,�l�.t����C�]����6�?�>Ss����a�s�������ɘ�����scw2�M�[��6^nn-��jh�C��K�6%�m�	��)Ry�}PON���j|bˎ7�[�fBʰ�D6�0�}�Tk�q�zA������_���n��H�⅊R\��7�z�m�^DPv1��~�A�zUZ�����g�k.&���J/:O+ז��MT����Y~�k����2���u��ef�~�-�k�o��)����8� 0 Sa4O[��j��[�C��cY�r��*����_6Vu��N����DE������
_�:[0 x:ţݝ���9u��.�1c����c#�1B:��e�'ޮ��ƙ���$е��+����^���:��Z��O0 �-��`c-���u��[��#���2�w�N�_z�>����sg�b�<�����Í;�����&,�9����
1Wa3C�X\���_�}��a�Dv�^|��>|2c�B����F]�rN��Q�F6�&�\m�k� L�y*>���爇W���y�xд�W�K��!�6����m�:���z8}#�����3D�e]�y��]oSe� �
��7���of=`���۾���G�
*�OcQ?�Ԝ����1��P�C�������X`�P�bP�^RIX����U�qG+ Ъ�t��VgV$���	~=���L�"�O�8��4�IOd'e	�U��;��W激r�w��Z�m��aI�?��"T7:6�J���VJ.�!Έ�pc����9��P�P��H�$��-������cJ/��O�FR4K�:����������J����c���b9B�:����J��I��n:V�#��f0�X2�8��w~'f[��'5Z�r�������/uyZ�����[B���YO�cI8����$���p��.A��)Yu���K��	9��aڏ�z��K�����7��d��P6+�)�\Ģ ��.���*��9��Mm\=KB�����\6߆�;����;;OG�9Y���Z<��ψ����}��u���p�����E`^=W%�|�����,�ڈ'�%v����̳?��'=n����/�r��م�Bi;��i0&$�ѱͤ"�C���