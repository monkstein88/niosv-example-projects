��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��0Ǟ���:�i�2����F��Cp�٧�%�VU��^�}���wWN#�|h2+2D7�ҸQ!��,�\n'����J?7?'��;�;��^�r��A�9h~d�2CI[\Y���T�Ū�	LDO����g��C��򤆤gE�y��l�'Ɂuu�4us����2��jC�^��|�7����(-G\=�=��dgR�|����&w��Vo����<izuk�<�~V��9�Nq�D��c_q!V��\�s�[�<7(X�Z�=�7~]�
j�x�M���؁ߎ��d dI�sry��syq�����O��~�y�?��=7�b�s'
n:���Coz����|���Y#>��Y��KC�gOYE, #��U`�>���&i��~+���l�&)9m���)"�v~�n�B��T�3�(k������QY�D�l�x����_<������y*f�o#�a��cd����V6�;/56[
��YM�Q��w�.;�o�U �o �l�B��v�^;�����*؄�*
''�f��]�m9��y��yJP��V�L�m���̚9�hF�)`h�g����>ùj���ǙB@���+0�dX�]j��j'������M.�E�8\_�p���]�-�-�jg��k���,/Kc�m_t�!�R����,3׺�עq��S0���|��a��ba}x���"�2YH��ct���L�M��d��(	u������mC����}�d��k	��n~)4�X3!C!��?	c�����ujݐp��g����CL�<ǭ�b{�Z�����2�m�.��̙�|A��}�v @!�&ӌ5h�P�M|�����"o(�U�Ԓ��,��Y�nJh�l*#J�N�hs�6�-�N�؆?K��ܰ�?>��[9����[u�CFS�Z������]�~�+��\��(�(�P���������:�i%ϥ^��KUP�Z?Lj�J�2�9Xc�T���R���5���^��S�N�6wF*�o����ޔ�jY�u�vJqPe��4ș��?@�sc��Rх�-�ROF4�p
����к]�5����E���\_�6zj4�3��<H��#�3�	����Q[[��X~�,�
5]����->j��j�?�vz�iÔ��e�A57;S|k�+<��*S��,�����R�����y�p]��IM�}��JհP7}~n�*'������4ؑ�,�1���ɑ[�3�
DD���U�V=�x.'I?Ŕ�F�Ӏlq���֓���tN����w����I���0ORStZ����<$�_�� G�F���K��`���4��3�`� n�[X^������~gՌ�C�Q��ܗ��.X{}g��$b4w�(Q��E ���*�j�ne'��/�Bɽ�=���TgA�a��j��0Ԡ��:h_Y��������V�s������607D�n��$�d��Ǫ�EK���
��C�e"*.�W[C#:�����P�����7Ұ�sm
�[�p���[��c�P��%qq��`"s�S�O�&���f<�n|tD��E�C�VR`�x8_�3��Ih�T����JgkbI֪������j�D��j骋�4P?�Ǒ�ey��q����";`�X�{��oԓ�,We�E.-	��gT����fMx�1V}��?�p<�Q��rn�N�a�fW��@�ډZ��ގ?���2ㄗea�+ԻSI�n�'y=�HP�Hc��'�0PJW�||Oӽ&�Fe��[$~��c1������*W�J@�X5M�PP�--�/�^��	����ﾧ�h�/��̽�<���{�f2#�"ͺz�5K�����Z�����(�GMiN7�#	��Uf�uTURR�.�k���-��dRI�ڳ���8��{9ZR�q!�2w�p��k��K}Ǚ�ķ��qu�(�y$B�ZPH�DE�����]#��M	#�&tad>S�`�O7gGC0�p)��66�wѰzۜ�]��R='遭=��i�=� �#\r�ňPw�5���R
z$�R�Y�+��{�Ś}�1�wɷNSt���t��?��C��{4F�ߕ�#��"�oM�:�Js��-�xY�#���=��M���CVZ��9�e閔"w:���Y�?��A.ӆ����L�P���Yi��.i;Q)�g������Gd2i��IGL�%��"�p��e�)��i(ó��[���	����I�fcX�>#Jm��B��_�5�*м����L��m÷�dj# ���`���
���u�kM���esx�ODU��-� �(e�����&����E�T�]ׅ���ʿÜx�a�����2W�:����H*��F�����$��*���g{��9�֗��K��D�l}�W���8e�����u�֗|���
T f!�:5#4�m�v5ʰS_4.�o�q�X�p��v�žW����!�n��p�J#��	2"�T����L��C7��3'� +f��g1MN�D��pw5�`9X\����<5]�����L�|G�H��z��RgBj��)K�o̖*I��?����q�.�؇
���@'�r��� �#-�nG��?h?��h�V~�)v;�ɍ*Q^?]��`G�G?�̪9Qk���7��䀹W�#�	�]��j�f �6��L飢q�s���#ȿ|��	7L��;�I,�%!�mDic��=/�3�Yx��(ޅ C��7%�F���B��!���`����;��?Y��8�:�ݞg`��h����P�>r�ak��p�i�����)��t(Mz=q&x�E��
.��6O�����!��� ��BxBLg���,��I����"�Qb��Vσ��b*\�U�f=���U��[0E�C�)X� �@�~c����b����t�\���r7��X���u�ܟ��L9!Q<��C&�쒐.!�\�b����C��P���������	^��N4�l@�i��v�	�ku<(gvtk���"n*Bt��Z%���[����j=�_AFns��A�F6h�����=������y1��'d�f��h-KT^�N�^�S�%8�H�b���e���CëV�2���#�Pqcd7ziL�q���'($�J=d�=j��S�3�d�+��ﻰ=���b.FAkg�d?�!)�rF�,ZN��&�K���(�iY�����m�O��W8���j��35�ݻ��9�n�¦�l2K�3,����bI�-�_
v[���0�d��Ϻ�Ci�~<���i�
,��3FR 8�wJ�T�n�;X����d���r�c#iM��$��鬽"}�ٳ� z�ڊ������߸��`��s�@���Çz��s-�Q^������q��0q��v�]�-_��N\�@�ԟ�i ��$,�}W���1�k5y�f	��g#�t��<<�@��d�J�:Z;�>l6j��X,�)�w͎
�fօf��1&z��P��E"��53H��s&\�|��9�+g�E�c��\�"��wP �[�l7l
���ey�n��x���
h�r�6�eA¸_��p^%�����t2�f�59��]i��!��)䚢o���ږYbx����w�g��1rD��z(/I;�@��!��� +���أ׼k��aQ�}��L�:��Q��D�/V6����:�����<��3i%-7��3�D�DU��Ț6�������;�Rk���Uq�2z�E���F��i
9B�E�.
_�a�Y,0[�qr�c���\gY��c��0�R�C��g��Q�f�����+�rj)M[X�xv�����X�V��~����2|J¿xэg�np�g
%�IGt�NxU+���q
	Y;��A�dS��X�}G�H����^XA��yf��U�W�q"He�v��)�§'[�����ƽAENվ�-�v�X��{c���/�^��ܓ��2�-������/��N�L-S���U���0�3��"�q��ݪ,��q��X�X�ǜ&��+_F2��B��Z�[+�?��S���{]P���v�_+�����&S��
���nh� Kk�m�=\@��+�:��tJp���7l��,X+0tl&���<��c�:�76gL(�nB�yC�ؽ�>��oˣf(K�_�>��uN� sǺP���=U���[O�&F�`/qO�Te�9�?��J�T[��\=͐�����p?���8/����c����"ƛ� ��h�]�*#��N)���1�������x���`%����s�ݾ&������M#�1$�w)��hN�>8N�0�a.