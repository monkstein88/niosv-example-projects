��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a���|�5��i�	F6J-I`�|����s�%# ^y��)�C{�)LQcf��Ae���k4��f���~���>V^nm�1��%�f<�5�r4�F�xdn�iw�8f�E�->7��J��Y�����#p���-�[���6E)zj P�_+Id�o�B�DCM�A��[vu�B\*�I���T�Ӂ�o� @�Cݱq�>��+W0�-�!Yb��I�zҭ�[��B�Iqha}Xz3o�����`���\��4���>��iB��G*��U<m�J_Ī�(�a��U,ؖU��U7.3��B�KdZ���b�T%�QU� r��^��;��Iы/b�㳷ag@��E9��7qP�]�� ���°U��q�;��~���҃F)-�(��P�b]�b�Rp�[��*�JJ�4��U���iBw���&�����U�e�*�NptA�[$,'o<*f,����r��&�3HBM��8�zSSX"�iu{�ć붲���o��p�>���A����/��_]~��{IBO�<<�V�6g���1�D�j�s���Q�ܾ�p�%��� n�I�QY��&��mEo~�*���&�W��ǫُ̊�K�8q)�U�B��ٚkҍ�������[�8j����)����5 �g�= ��Ui�R!:g6�O�����o:��ꚽl�K-r�����;ƗA���. T�-����7:����_�:7FxZ�CKl�Y����
9��O�j�$l_r�RZ�s|�TW��FKFSa�tL��p�w�_Vx��b��3���U�Uv��T�'�WrD	�
q'-`�w�n�un?f�^&��H2$/�i�N�+h5S�	�(�Ύ����_��}XC&�5����tț�pā��8Ԧ��P�H	��6 7�J�"�����ߪ\�4��5։WA�ؽ�az���jL��eTz����D�Lȝ4b�5�����3V�Awt�z�*CҖ�)�����l�v+x�����W m��.��7w\+���l�GU�������G�9��e�@t	�>7S^*fɥ��U��-H?���qE�>_j�*��~t�VJR{��#���-��$I�h���~�',s�~i�|�"���'q�
rZ�8��&����%W j��dtn��g62Ϧ�����c�O��WY>�h4���''q'�5R�A���1��O����u�*6T�rx�*[���|�s���,o8[V,���9#qv�k�ڗx��F�ͮs��B���y֗�8�C���
��!M���lI���F��E��Sw뻲��c���!���� �NwB*ҝU���H�։��`b#^�oQ1%��z��b���I�����C���v���@����ieoZ���0Ԋ�["���/8�5�f��NZ���oN��X�@�B>1��=��s�uh�7�<�0��Q�����$~ )�[O�����
�-~'$�]�@H�yGE�&�HrfM�-zC�eӪ��M�.o����1n�f�*�� >_�8�j�,���}�ϝ�㥣w��d�G��7cNPu���ӳ��]���;6RK]'w����n�d��3΅�|���b�~ģ�/���7v�zWۑpd��U���2<�/�U^����Tmƥ�4Dr��$�h��,��=����Od�1��xD�)̛�����"C�l�I]��40�ؾ�g�F.9�^�wz�>V@9-�}Oأ8N�0r>**B�+��)��̬�{��=X$��;�,Ʒ�;�cU��|G�ʝ�4��V�ɗ����BL��T��0窈�7.*r�F��$�:Fي�AN6�D��C����+	S,���Y2��L�̈Tx}�DP��x�D�Z!uE+��y���d�qh0x�7"��<e�������ȍ`�P�z|�BH#���QU:����L��<��3Q��[�Ըgli+u��5ђq�۬�O���%4�����6�Q��Z�a=����)/v����,@���� �[G\�2A�J� ��W�a���5ئ��N��Q�ÐۢE�4���~�7m�2U�N�Jbh�x
�x�!`�|��Y�`�KV����6���^zm�E&a�Q~Y[�⽵l)ċ���R���Md���mwfF),r{[�%��v4c-U���,��K�C�>y7� W�҅KJ�ڶ2Opx�ߒ��s(P<�:�2Í�#di�W;�(̜'}��m)����O̘�K�s<y�s?������>���\��7��=���z��j�	1b="���t���("���md���r�j�-��^H�bxe�b�%�^sR�e㭠؊ȱ��Dp�e�I�H�uU�R���!���ڱ��L�J85׌��	�]�SዅQ�h���9�<�������`�L��l�_�<��I���Ĭ�%~����r�D
���ei�#�)��z50,�̈�  Z�a�����aأ�S'%c��m��v�p5VcD����jŤ�[�u �@,54l��5��������c#jE<���������:Ā��������Lb|}Qx�m�a���T�e��z7��Ic;f���#̳ �e.WW���v��Ѿz�ӁCRUFG�y� ���yr���A�{3�I Ѷ�}�ƫ�I��c���
�M��gY��og��I��c�]^���+s�	5��)�
U���|bJN��965�����<hs�R�D��u'Њ+���}1���τq<�nG�5�,s���)́����'D�uë�7�E�s.��������}���e>����J�_ݎ�/zl+#�M5/����%�yd�2ۼj�ZM��/ʕ��ft�
 ��Į��i�};���'�<F>��u�ɵ���Z��%���͈>DA��c��4�SC�ݭ3m��D��]�^���%��J��Wv�� |�MX�z'ǟ�Iw�ϛt�@���qt��]f=�(z�Pz\
TU�[�E�f��fa<7i�+�Qĕx�O�/lh��D�!|���؈
�	�L�ZLԽEN���o�>s4��ف%�z;�%l�����r~f%A,.�@b>�Dk��A)�9���Qx��HT&FOj�eBl�5�Nv��N4��Ȇg���z.jO"#���i�K��5�C�\X�������<%c�dܮ��$��ô���5��D~���4�=(�Mmmr�+�!d"s����Aȹ>2�Q������Q���~�g^w {���ǟ���Τ)6��64|����%'���8Jg4K��2��D���N.��Y��q� F�ORU�,ȥ��M_/��X�����xR@��B�F5i( ��|{��k��2xHu��"�՝���4�H�̠A�G�R<\H����6e�O�}
�4���:Ţ���T��Eզ�]}�'��j&'��EEg(a��h��{��dK�����Y>_�#��猉�d�X��kCΐU�[k[��GDd��ro�v��5�^3��S��P8�iZq��2W��V��_��rl�"l���7�VU�=���8�<�"��B�j�_�4P�x�Ez*E��E ��9�ی�������(.G��`@tW_��K-v;�,	��ֵH;>j�P���n�P7��G�Q��T����Fy��0����w�Cb?�1O�Y�~{Qj�T�6Th�Z�`3��ܬ��"Rw-y&�"�<O�<��ԋ�n�����F��7/������Au����x��Z���m�bA�~*�;���o�^y�؊���T�Pk�'�* n�|�l���@$�K�Maꋢv6H�9�t��t���{�؅�/�b�/ ��=���X�G=Z�F~[rm�O{���Ɩ
��XOI�4��Oձ �ϓ6��aE�]�o����+{x�y���4�-.������&v4_�}?�M?��H:Z��^uw1��\
N�N�Cb�V6�ލ����8|m�p�̌Q��N��+�n72���f�a�UGRΊ?���ۘ0�ZV@�m��
�d���ܛ�k�U~	���kV�_�ѽKY:�����:kT7LT�'�����}k�/@+�e`żv��˩+�?��g�����>��O���z�:m�Ayb�h���u3�6�p~+��!�Qdv�`��O�HK�'S�>@_3�K�?ȾE�[���k�Å|�g���t~��;o�.���#�>�j&���C�� R�f����\�De1�pA�v�j@�}�����QD���ы3W�������B�OE<�^b t	�ɿ���|Ļ�6[2]��-=p�Q�L�����ȽzCNm��	�������p\����wx���Z�}�q�~I�~�Y��5�]��$-�]r��+p�411��:
{%�(�+�K'�FU�o���w_�p�c�άKM"��#2\��NrlA|,ؤT�8��g�Cf�l$��(s�jV���v@�%O���#r99l�"h=9���רgfힸ��f�4k�:��ly�.��Y�@�x	L-2��A5G���x=��OǕ��A��&�ù
��F�����ZWO���BY#xL֩���p/�5X