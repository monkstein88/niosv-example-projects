��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a�����/�	v�+����@ɧ-3�����Iz�t�܀Le'H>	6"�U{��9�bEɤ6-�!�V��s� ���m�|����~μn���}�iԹ*VC�4���m7���-� �7�o�d�0wUQ�z:F��:�����wq9NI�|�'����b�C��Ӥ�I��Cz��,�7Xmf7D��3Y?&L3�?j��h��o�dƛ�0��H��A�H'Fp؍TCP����W��p�/MBq��� ��,�NG��Ӣ��:�6K9R�d��Hf��o ���]��0/���Q�'�FȨ)��V7Ⱥ̀;"ݰ����g�,I=��^?i�S�@)�h��P��4��+���'� )|<v��$�i,�)����Tw����~A,�i��Z�lput�?>��U���T�)"R���F��	&j�M7����G��~�?B��\���jj2�#WK;������!���]_�ڇ������`gF ��jΥd���HrG�
ܶ��?xX�,0�Ֆ�'MĻ?���} ��X�@�o��l$F,�)�IOqV\ݨԯ2y�Nȫ�D�>^�XE���VQaCp������a�~7��Zbu���/�cB�h�3Y��Yw����VO �/C+2kT*J!8-��?\�N���X(�?c	S���5R��P��m�R�´����ʚ�&e0�G�x�d��&�ZcfN8YjQ�!��K�iW1�s ��¶�pT�dв�t,�&��䫓d�Z�`v`���V�qFE�T��E�·\��� ���`��1�`�b a�D�.��;�����VBsC�"4��:gƔ�Qт�I"UR"`��҂/��T͠� q@_)���A�Dh��qG���U,<�	h��v�0y[FzJRH��,�Z��kā| ����Kp�/q��B�N1Kd��}r�U:�Cb~�P3�R��o�h�+!Ӓgb�S�0�ήSg� �^V�}r���T,�V�t&��y'��Մ��T�l�ڡڻ�H2���<���ˁ��2Clw	�����?�p��Fw�9R/�LY4��Ʀ��z�M����`I�9�:�ELn����Q��ۥ����J�Q���r�[�S�S���M��<N*#��5�}+_��M��ؚ��|�5\H��VPe��ِ�x��@/L���5���sl����`�#�jS
eѐ�<N�gR��A�e�y	,�A��%���+dg8�ο�F��&�gޜ��;
b��� q>N����m���<A�ϔ���5��q%�B��7q��1�{��?��a#4�8Fԥ���I�y�x��J�k�''�.a%+5��q�m��ny�ۗ�p,<2MWc�Y3�K0� 
���}!M@�.���'߳B�vd���ù�ю�@�{�Q�\�0���4�rw�А`�� �b������/�T��m�Yr�H��������S�67@T���<=����#�oŠt[�k[��.��3P�h\��������!�Һ��(����U����o��~18z��!E�$��X���{c���2av.0ǌC���8��}�M^����\�UӰ3�咞��p�H�@S�W��
�F
�К�N����;3��P�����&Ѫ��$�n���m�\����{�)5�H$��S�gx5�$>l��Hx�n �~���R�Lt��m��>�x�(W�͉�HQї�@�PZ�P��F|���\k���8(W^������&��-@��AT��	��P���W���mKL�4W_Y������
�΃����|�Gb�勶�����7Bc�̳���XEr�/��&Y
]s��3���s��>��#�/S�����O���;�ܛ��b����w<G�&HҪB� b��/��>��f��2�Hȍ϶u^i�x�&���
ݘ��&���u��J�[c���)��Ή�A��l�m+�M�7h���/�0����^��9OKs_-���}f��kOjh4�0���vm�'_��Y���/Lf�f�`z��V�\�՗T�ۓ}F;Ѵ�3k�1��+���E���5�_NA��l�;���Z"+��E�3��I���eȿ#K踬W1�	����u'���HP�E!�ٺ��i���E�Ѵ��P��~��z�CR��"�,���sڟ���ԊQ� 2��)�![���!��m�`T���~��*`�C��In����˗X��ti�b-��|��������z�lt�^h\W�Y�lFD.�d�y��b��Q����a����N�ٶ7h!MmY/V�J��zދ�3Zm ����%��} R �fŭ�.����<AO�����r��������ԋ�;415L}Qcx�U�#$]
ǽVq�Ԛ��Q}�|�B2|��Xh݇L�ɠE���4Z�f�Ҧ���lq�*fUN�%��(�����y����`>x��ȩ�q��;L��G=/��jׯ�C�Zc��]Y�w8�cn�z��z^]azN6B�K��M<�M�4:;�'�dJE�j�Na(bF�@��*����D����o:������l-åO����<��E~�/�JC�;2u.�)�V$�Ѐ�`���r9�O� d񄜯a��|�b+;N�mC!ߕu=�<�6б���Tf�T��
Y��}�#ze����������%6I*.�~� �A��OǢ�����V��͍+�"��Pu��"zFj3�7��O�ZU�~����2���)=i~�Y��f�y���-}hW�>���\�$��5��wQ>'\�g���CX9�<��ܜC�"�a���D)��G��mz͆��!H���u�n|��������Sk&��4��*�ƚ���o܄c���b����i �O�U3I�>��)���w����C������b�$\7b�D�����Y��y���:�;N����/p��R=�k]	O������
/�����M�-`ͫr�~����P��~�(���K��K�L��b23��+�ߜǅƩ��}�g&`m�LȰ�^�1����'�2R�4�
�0���(
���ȉk��=���]t�\h�N��[-�	��_ԂZ��#�]l@�q�C���R����)��W�A&���!J��.��x��q�OЧ��V�b�y+�ՍX���������w�BT�~����]�P?c�FwT
�hj����c=��4o����z��^5�g�ϴ��1�ŭ���Ǎ�t��W����jbD�KC�{;��,�Z供��w�c���m�= YN�9�56M�>?��xI���ϐ����W�G�qv@,�;��� n�Ξi;7m��ĭ��Op������Un���ɤN���$���-y^t�X�2���{[�fwA��5w V\#�	�G�m��E��v� �SQBX+R�c��8Id���F�Ma�&�3��*����b¦� ��t!��P�{63t��}O�y�OUZ�j���^e�6AQaR��Op/�:�"q1��1Unj��H�p�:�/1w��P�Uf��u-�C�TЕ�/����<Å�W�l&oi�3�N��b�Z=�ea@J��iS��|�a��+��5O�R ���xdL��R|Z�&XH>s�ose�-P�6G���b�{�K�P��C���[l���>��]�C���řE�L;��
���GkaYg����������|���º�B
rB�^�!���[���3�ű�s~.���͹툸N�#˚�st/伽b4n.�]yus���x�5ۃ�q����Q���AYsQ��`4P�K<@jS6~�u��\��2ɱ!���v�/��a�������ǅ��qgǓ�Jn���I��Y���9�����8�Y�\G�n���>n�]�f�L���uz�i�S�a$c ��JUp��t�+�|7l���Ƌx^���B��rh��(#c ��F	��=�k��)޴��2���� �o��u��S$Z1�;t�#"`��L���E5�iI��+�l?�m긃Z� �M%p�����K��&�>N��f�S0W���S�ٔ>��G2������{��\pw����PI� JUV,�fr!IF�h w�{�=I�S}!#D�&��\�'%|�:0���vt�j�ε�;�K���36V�a��uZ�[�>F.`�T W	�w�]	��b[5o���v ��ՙ]a�G�+�G�>�
�=�PIVrn�D42p��!���c��Y��������o���PHt�VK���jK��#�@�}-qd�;����L\r�����I.���g�\Q�֘[p�N<Ey���cHҼ��I��Vo5��/O�a�(p+��s�nGT�̶��9�w���3�y�&1AHު��pHJ��K~ޒ�
����3Dt�$a�߿�9�,��R��B���%���잛�M����\�Y΂���u�p���+xr �(%fO|w�x��P�����O�߉4��<B9eTY�w��4})�����f�`l�yO�����[�r]XfɐN[%>rf��,6!n��B�^m�|�������716��alK���� ���|�2��}�/�9$K�f��~Ji�Z�����Ϧ�x^w��:�!]�ߵ��f��M8�]V�2�c�+�;�lO��m$I�k��g͛vTZ'*�EIh��0�$b�^a���hE�T4g����ԁ��uB-�~ޔ��0��G�fJ�������G��`���OY�ya[� �Ug��*�ņ��Ø��
��?���������B��ϊ�)�;�vp,\�@���� =��%�Fzg����־��@r
��n�_�OqŊ�ݰ2���Qi� W����x���΁E��n.h�gu��|B_)e���#g9~º=]3�z<�y�J�(���2Gt{[v�����\k��gl��Hl�+�ߢ����ͱ��G	́�W��re��b����*Y�;�i����J �L��D�}���i�}9�j��af����x�OJ���0�F�6b���ԇ;��Wr},��#����2�l�;���M����no󣲴��y@S�9E����.f�5 H&��~�ц�I<�m̌0/N�փ�7��	��;�svd����F���%�T `���鯊w�Ai[:c�W&ÐY*"q��X ��q%�_Z@U�϶K�WK�bW�a�rۓi��ҁ화�z�[*�RK�zߝ�� �mF&���G���u��^�������1�U�Mbn��R����W̱�&�������d��5#P�aV�����{��rE�aŕ�g6H$G��7*�tC.n;j���X�H1=i6hA頴;W.����%�۬���k��[[Ь�УK,����@r}d��s!+�zG��L�������nso;���5�6L<�C���K)5��lj8�Av<6F��Z��=+��b��ҫV�p��-|:cD��I����b;_�	i&@ ��\�c�N����c>�%G���$�O]JOfJ�(� �����t�>��^�����g�R�[!�������[N��w��qCP9�w��� �F�yȢ�ah��!8g��_]�+�s�j��b��fQj}*��M[���1�&�#��巌Z�Z�M��Tr��J��~�|E�F�.$����֓��p�b��G4�9:����c�e\������4��uR�V����©��z���̷�����������:;��+�oVEтv�*n��2�)�8=S�$�4;�f�~:U��:aA73�{6	TkVj�@��O	OխיV��c']�k�����3ce�3a� ��Ɗ��Aڊm��t6��S�CVt%ǶX�J�}�� �椝�Z���"�Ʉ�kOd-�"��7Iy��mK��"������d�u�Jp���\k)Di�A'� �p��V���8���%#��/o^����ç��E�A�h��0�`8�i�gf�:KX/7�j��Hf=xJ�q;�љ�ƨ�_����w����&�����"�/�s�����	b��ܰ������sJ=���޵T�^���b������q�׸� � ��hMPa���@?1�ϰ��,ǎQh��/��"�%�k�C�Y`�s�`/Cm7�Dj�󅎸�V	�u2J�Xx�MN��fys���H�ͨ��$�@������8�=޼- �ރ�,��4�XƠ�-#�Bs���Y	��[:�}�̲�GZy��X�Y����o��c&����L�
�y4��6��� ڪ� f-Y���?���r�����C�3�~fZS�ǟw� .��P�E.��s���g�����XS�g��n��Ϯ*/{c�L��O�@$:땝�>o<֢o�hSw��,F��w���h���in��d��[ƖB�@�:�ki�wU������������P�Qρ�`n:\��#�G��<דS�c�����ϛf�/}�a#����X�n�j?����l��>ͅk�.`��{��Gs�7��|����Og0���7������ �L����V���OG>.Q&!��α7v�6��#��,k��1�Et�#��e�|��VJ��Pw� e�˱�X<��&tZ�	f@H�C}m�Q�.��5���l�
WC6��!J��}��k0�h�DE,�#�<2͑Ó�:�t\XTw�BL>/��� 4��������������P`��-����.�Xg�P�6�= ZS���b�ۚ�?q���z��Dw�.�M��	�ǫ����
�/��Z��u;fʑ�BЇo62�3�KM��[d��v��U3�v��9��>��W��G�)�"���; �)��Ok� ���1]�	�G��¸ҷ~';�+�x[�+1�o���� ��E�7��T!�t����a/w��zV���$6S�&�qu�n=	qӺ��� t��5�K0&�G��5B�JN�6���<g���d�d�!!�͌e�ʓXU7)B��N��ݵ`bO�5J�n�w:pz�| z�1
�ϳ�P���~V] &$)UT�KT_0Nχ�����=ӥ��MZh��*b��o�>�y����c}l��<t
4{V�%`�¹LNV�7'��� �0�w44���]x����Dʬ�0�~ǶW�准�| ���g�dJ@���\�P���e`�OLӃ��*@�9�v��cH��uM�'���$S���&Yث\8d��+u����3mv��˒�2��r�_���������������9[�Y�J�pi�����7:��+Cc�^��Ք� ��F��9�B��J���pu���V�KA�d�iNO{'�K�]�٪[#-�A��lK��xT���7p��rHN�\��v���Ț�惹����?��)��ۙ�4ޭ|�S֕��D	>1P-�#l*`#�
SJ��yzu����a�T���1>�w���Os	4%�5�Fr�FR��,�R�Y����b��4	$�<�Œ�X��P*X�n��_�6�]q<�x�(Wt~h����I��(gצ� ʧ���kL�Ϋ�W(�Ha���p/�
!�=X~���&����xz�S��_nMӠ��.H��Tdf��]fi�X�pT5��)��QJ���DۯŪ܅,�L�I@��B��cI��i�s���&Bs+�qt}3w��Pg0-�8���4A�N im�� ɭ�~�.�[�2.�Ua�F_`b�ð��de���B0�3��v�������4���M�����[}�߉T@���q�*��% )���j)�Q���߼��f������e��D�2^���/�ư�\p@D6zI-w�J��������M�$�5Sa��V*�:1l��b��r@R*��gV&���,^
�.6����&r"�T�(K9�.i��7��ͥA�NK{+���ܖũ�(�m��(=��,t����3�]�A���G^4#�����d����J�qc���!t�Z}�K����l�P�Н� �?"H:%��@h�b�-�k���a���.JE���GeR8��\#.��"��������7�+'Fn��<�H�X��K�$`�
�h���Q|��������]R�.}�^�jp�u�h$hD�@5���︤x(�JZJԜ����9K��f8i�){�(>�n[C����)j��n�1����?ie�(����>����Ѯ{��ps�.w90���L�<!�R�ts�f����{	�W֣�Ke��2�����a�>�M�ۭ������Am8.o�#��FxF��4*��SQ��(�X=-��9�\�I���6�j/��	r�D�<�4\�5g"�Y��I#Ĵ���Jc_ǻD��b��\i~y����w�VF�s&�����Ex�4}��G�3�B�*��+��s��c,i=|M�ع�[O�� �H�Q�'_���JU�x#���7��N��G�]� �ha�:@�z�w���Z+ֽ$@L���g��×w)s]��M9lg�,-�+O؊h�*OG� �>4Q��D���%l�U�(�oR���vԢ�:�x<ދ$L��I����p�hx�O�����-#"�� ��{G�b"|����RMmcB �&~Wb�6�?�rr�`�-:$c��MN�6R�be�d/�7��h�u�7�p�2��j�d� -!�e�i_�	:)�9UU��	��F�0>��LB	��#90�5�WZ�x�i�^�B2F���-�n�QbL��-��w�f��Lv ��4�l�����ߒ���/<�����CN���HX2�Z�����	�c�I�.��T47^�h6�֒/9�� ���|@2����qR9�.<�1�F��Y5;*����2h�,s��k����[p=���9%��l��H9t,c.dk�3=Z�>Sڧ�2�.��A3�Kq[	��|�JR;�y�}E��Oj�<`=æ��:��G�e,Z�쫸0�H�t^��Q�"2���3*k6M�?�-�����BZ�`��i�	�ar���=���]g=EDB�
���q8Q�/�����4U߳�ZD����S� ��{��R��2! ܫs���5��H?v����$B��1}m���r�3;�L4M�6��c#����^v��h��+�z;'�g�S�i�!|Dn�B7k*���;���: .W��]<fT�y���������i�|ne[�ys���ĀV��K����R���=��mYXCD�bĸv��M�-��(&eJ0��lVZ���ә�槬Փ�qJڝ�f�3'Q������uo���@����'g�<_�G5����� �&:�{��y@��i�8eq:�C/�����BQ�K���XVK���W��r Ԑv'c��[]CB.v*}0�5���u8�wQ�h��`�� P"�����f��'��UG�GM/�u`G��LW^�Ջ]��U�/�0*`�C�(Y""�o�EF����,��~�־̽>��"Q�<��H'��5&���|�F#s��"�q���ŰD��hg'���|�q�2EM�1�x����y}��\��+2D����Lٱx���h<�$���Wz��P�aKZ���h.����Hc���c���pX�������� %�x��u�����w����1G�TŶ?�U�d���T$ƺ��Z�N���z���NWq\�b��/šsD��B /�*\��T�
�t~b�N����P��$�:z<&wk������
�1oj�?WX���s�_R
�f��w�P��Ǝu ��kK�dg@!yи����늋��v����H�ov�ӃUt���O$]�����Ǖ���/�Ĭ����u�pcj����EԀS��^�O��`�x��~�6�
�	KX+����[�ٿ����<`���(�Q�q��i6xJIcp#�����?0��S�� ��r�l����i��E��6%��\���V���@Vsȏe�'�Gd��>��ڍ�td�Ip����H)��ZL�A��
�Aķ�O�u���g����h kL����EV�{8�5����p����~�|6�㐇�Z�Ӑ�T���x�W��)W�\�"BY���u�eDUQx���4Mp ��al�BaI?���y��.��D�S��ė���d�>�O�H���\����F	D�������a�-?�"��;��0��v�f�?u"�^\���e������VDdG�;�G�P��D�6��8j}i`�e�Xd������p�#8���k����7��i�"Ř,�>�j�#`��KRB�A�p������?�����d�+
ANv�DI�����s�L9r�m4ΥYC��ע��0���g1�_�1$�dQ0�Ch���
�O�y�;m,:��.1c��K�����4�@Ry�tԗ��la ��c�X~��20O�ך��-b$��P�� r/�2k���u��K"!�����)c��Y�0�L�m*����"�.VG��+�������T��]Ͼ�I��,�+Sȱ�0���ځ�F|��V�x�G��1��z/4�=��K��[Ѕ��|7�l�J5���5�Z��/��!�j�;��#G��aaŻ�p>��=�a��Gy����ݩ�b��9�`�m�����7Ѽ��|�4`/>���J�!8,~謷�	&>�Z����d��p��B
"�/(.ۙ�=��*�JNʹ�ej�0�,&���o�zNi�u��a�e37�mJ�!���х�$��*�8���E�#��Df%�z_�j=��v�bVk/����H��4L^����E� �=[I���B�i^^�bTkAD�f�}����mU�#)+�8�)9V��1�+n����<5�ZN��	����d�c��nA"����z�l��њ9ϰb�ܪ�b޾�1 �l���w�\$:K;ed���8�Ԃ�M�ʚa`Hݸgrb�_\�"1:wp��I��s�����|�AB*O� �����֥+${���w���~��Gg���бUw3x?��aﺽ�|�X����6���~����s�6W�IB�H����\�3�6Q��D�h��uɐ?�*�R�x�S(�E9��=����le��n-&������pUvE,Tn�hu�2@u-�D�x��~h�9#13!_��_��� ��|X)�
旚�c�~�,��(�M�q(�y~�U��Gl4�F4�(/��������K[���Y�ԑ�5�/�F��8�\5�ʜ~���^�2�S��S��+�Q��`�o"Kh�jcX].Ĉ�C��U�kN*�^w�,�a>4�`��Yqc̝�T��߿��ݝ��@�	ɛ�s#��)�On;�J�q�u$��M���p���6�F!_tC��˨aO���`����wM�v����y�y���YdH�><��9Yr�x�F�9w�@���
2�!��Ħ̓��_�%�n����m�-o�X��.�[<���w1��
��HJ�!+C/�����}����p�Q�f��p_Y�ŤB�Z�4"S_0m�
��h#b�P4�oC!E7�K����!A�CŬ�P|	�+ �{���4ї�G$�֞W{S�ϰD2���=f8Y�C�������~Ue���D���������wJ�'�1o���x�aKV1�g���!Jx��S8t,����B��M�}��CǝY�4�Ry}���R��EK�,&��C��ұ�Wq/)�zՎ���wQ�ʗ#�n�Ǧ�ű����~�r�*�1��ۓya�V�8���7�j��x�LcUTʮ���B�ή�z��M�*g��#��	�mBh�댬���f�:�s2�e�?�������.�&yAc#T�6�1���֦���ms�-PO�W��^w�كv��?��B�4�!W]C!�}#)�X����|���N�S5~��P���3�|S�cB*�R�&a�M��LNu$��A=I	
��>��,����B@�,��z��f���y�z�/�'�n��k
��/���ő��#m��_��HϛE��N�ɤv>�ó����&�I&�O���C��`A�i3�HW3,��K
}Q�5id	ċ1}�,}3��xA��H�{G�S=��ؔ��{����2�J� cT��[��t�@�Am�t�[�6�<\�7q���s��o�/t�ޤ'a�5��L�Y/��Y�֔��"��$�L�W0�j�9�EW
��1�,M��3r��h�߫d���m�Ps�t���%�����v3 }b��8�聺Y�ߟoX�-���;�v @�k��Du�_7�5{P�8_Hg��՚l������UN��wO{�j����8��;���t���=⪺�C�ra��Z��e\0v�0xE����܌��-9�Z	O�;ٝ�Kc����،Aw�	4ߘ��� �",V�5�jˏ$����8Y��59��٨0Ɩ����z��,�|B�5�p;��.���Wڄ[��p�5�B�{��u�IwȂ��{�cA�8��\-�ڹD"��ӓ��٘��v�`@���|� �Z%@=���q�N�;�I�1��fY�#�	�xGyњsf�^�m����`0��8���oQ7�)�!����\f?�ſ1k��	+�_�/A�E���������3�e%��_��i�ϝbv�/-�HڽbyMd:|���_�.�)5�e�Lr���z��=y
��旃1�sW����S�osAnF����|��d=���X�D�<��෸~\�A���X�὎�t�+Up�Mq��n�j���:
AX@�[8C�I��0��͍)���`~4����2&o��Ȯ��ܢ+�l��Y�xV7Q�g/d�����'LB�;�=ܪ�Kx�PN��0�_���d���jH�	DfU���s�`�DW��&=^J)�.|(�/f�����ҎR�MD磘1���U����~�
�D|����=�B��Ӝ.Œ�S�ĠB�n����u?��߉B���V�1+����0ud�'�M�.|���P+������X��㵢�FݍH��{$RXD�J�T58U��0�x^����ef�5֦��K�2��,�L��1_e,f�&'v�S�u��h��R�<�|Uo>D��(��կDYo=����ĥ�~�8�;�cg�|�B�����9�U��ۆ���ʺ�
Ous�0��ԣ�j�'�P �- �k�v����/�� V
��/�2�>�>�V��`P��$����I�9Jʪ�˗�[�ҏ"�
��Z�����϶3���}��֜�-x����a@7��(�nqg/�����5�����;+�c��x��+ف!��� ��]`��%f�\��4�8���ŞT�:{U��iA;��>_e9�9��N�J��S1ʃ���H1���7������S�^l����U���}y�� +׃����dUT��~�)���9���|K�t�y2�};<�^!gP W|�ר���(w��D�PVH���OD&@��G�~�z��hB_ ��q����"�0&J��8Ҡ	x�%}�qq��E�s�P����Ht'Y�w����p�pF�W=�E�sڒ������9eKwg�6�D�.ޒ����)=�t����<r��*bj����Z�Y�Eﭞ�8�RM��Ԉ��K����8�����'�Xu����"�z�ɳIӳ̎�?Y�ǎ�`�x�������Ƴ�t/�|�&��˟� �ќ*Eݙ  �"\!���U���]l�a�ZW��>�k�s%�+<U)���ҟȩ�*c�1�*��9rH� "_����ّ2�ys�3�`d�lu��	�3�6��ۚC�!���E5�i�>�*"nI� ٝ~���p)V6W`V|R�VS���ȉ���ڞ��^�>�-�����
�+�*�`厉�g�i�A�k*Fz�:>6�Wg�|n�W������'�"��ip���j+���RZ�]g0� ʡ.,����݅Z�r=�d2g��$������Z�����k��.� �gFO�n]4r�� gVQ.��	O��ɪ�A~y	�^k%��sk�fgc��+M�Ź��K�7ou;: _��7knܰpr����Yca)�J�s�P/�Z����N0����?��4��ȫN`iT��o�z�bCo������<%-(�f�F�ѡ�Yi#<m��z0WH�0CƷx!�l7�f� �bMo1E��t�G��ww��)��FYܵ��V�.�t�S��[<�&,�u��g��+#U�m�>/��/��]��8����9���Vd�#��*�`����n�а�ct�|{L�u��zFQ�$WʜF����+s<�*�E�΄�Y_<fe�P(���k�u�T�+f�eBIp�H�r����5ͪC�zYq*+~ٯ,���n�(5���(�K�N�?��6����V>�X@gC��dHq&��^4����ɕ���v"��k���.�]�:�:f���@�\��sjb�� ��������r�s����e��+��Uw]ٛ���m�#�\\?��_vOi�vm$G�Ӥ��o�=���Ij�2Cͬ
�4�3�������E���H�IP��� ��ת���ڵ62�t�n�H������MC+�^l�m��n����O�W�Y�s;	i]����ؽ�z�jR�D�W����]��(�t��G�0�,Ԧ�-�`~e��ٌ�#�m��ָu\��i��fQ�C��L���Ǜ��J ��)8I����Ƅ��<�ؠ��A�:��U�W;1��t�yĢ�(��M�$�z�%�U�r���ɫ<eg��-�XA[��f��f�?˔KR���f��q��S�ଖ��Ї�$j����l��YZ���5"����U����`��5� %Y��:�3�1%��ƞY�*�զs�\��<Un9����#��V]1V8��Q�MB���|�tx��� �*B��[fw�ӭO���� ,��FdWu�����,⅙d��+�bd�,��H��'�Y��pԑ>h����Y;�d�!��Xa�~2m"�} Xg(�҆Q������}��T�a��sY��aӚU`-�}t�2��0�?
1���>���
�o%�]خ�h*Zx�cg:����h���66H�G;q�h���!g`x�z(����V�3JP�[��(
1;T�����<�2�>W��Q���X����ݓ��NLW�--{d�a��7�4���OFi���P0C�4�h#�@t��H����؆p[��6��Y y��ԃ���{|�᫮��Qb?t]�V�	ʔm�z���m_�y� �L�Eh��u|���������0���nG��O{�9�kB#�W��Ю�ϱl�!S�*{4͇�m�C���|�4��z��󸭭�G֍ ;vJ+���#�Y�g�`*Wۑc��S�b���9�Q�V`��>

.(�~ށ�L��M{T�F�K�s&C��«�[M�:�?J}%��fr��g�v���c1��n_v�$�J)y���j� _#�l��	�̬:�ߘ��`���s?]��ȡ�=��ħI���b�B��+7�n�Q���t��C3&�����.-�Q��ϼ�M�3��!xw�+�~e�-黣�\��LV�J��C�`�s������!������� [lw�����c���qN@�\V.(tn��9�f�@�MIJ�~��4��o��g�-��ΰTM[Z��Ej��#��˖�Y�z�2����0y'x�R=��x�ןqI��sW:�
�J�؁�e:�c�O�Qʂ�,<$�fA�������8��N̼���4���B�X,�@Ve�X�1�e��('' %ֶ��/4qe�ء9��p+�fۏ�@/�l�U�c�P�@�B��xM�C�1����T����r�-��+���00����`�O!f��ؾO!���4�ɔ�'�`�E�[�f�'T;B�{����D~E��ibM���	��',��bj/�i�H�y����ǽ�Ĩ	��m�؟��qK~��t1�D�o�7*\W�~M􅅥����� [���8I&��,����*��!�����S9*�*�����Z{0z/EÒ���%׌tl̠2H?�/~$�tYoS���9CG�~l���r�����K����g2�l [�<�=W�X�f��Lrr+��HʟyB�8%פݨ	^@3��0X,s��a^�J=eH9��FW�^�Ͱ�*�����w5���lkb頜i���ksg�B�
��7����g|�l�x-�S�:U2����U�s\�v&uuԙ�g>"��`�!
�t<���G���N�PW��g�(Y���IB���0�k@ɐ�υ���W�@@q��1�'�.�S�2o�$�p��c��bMV�^FN�sk�Q�i=A���:@�Փ��G��zˣ���^җ �����P��]�����{7�o�#��X4���T�3�dڻ��\���9X�̦��mAŽ�É�Csk|�����n,bX��h��wH�_�o�(G
����^�g0���An"@�E�FQ�K�����`?Z,)�_ދT_���� o�(ez�*Y�Ӌ�<i�B�g��wߙ5$�f=�M8Z��r��[�����[��n�yg��P�ʩ�K;�߭�]|d���
z���Ҥ����f�6Z6�a���#��x�v���(�.��Ʃ��ͪ�
П��`;h�Y	v+����%���W� ����[�
0ns�۞ѵ�ɵ]L�ɂ~cj)���K2�T	a�/�.Ä�����La��0b����<�1"d�̞��Đ�4��}�B:�K�������i߂X�&BF���������+�I�i���h���X=\�?�H��fV��Qe��w�+C��Ԩ���OnS��6��!�/c�,�ۑ5K��7K��)�}>�ylB1j�_�ֳ�@���IW��g���`U����+1 @ڹ����$�&�zj���4Ԁ��>4�z����vYSN7X�V5ײ��Kr� N���
��Lk0����$/*���Dœ�X����5W��U~��/��'iGDZ� ?�����
�W��S`�:?�Rq������BO�Z����S'��z9�{Ѭ�hsLΊc�����R���P�&��O�,��{��(���?H.�-��݇1��j+����R�����k׈-�g���ܻ��i�;�~���Kġ�R��#�����X�\v'��+:�S4S�����u}�^8�c������H�%Y�Ќ�:��u���J+�I���@�m�HW����@��Xf�v���P*�3/�ԋ{�qkx��"H��KU��O�#h:��QP��N���(x�kf!&�0��NlN�r�̝���,��%�9a^c®yxǣo�i�)�ɧ����o8��l��+!;������L�A��Ҕ�</(�|�z4#�q=�1�
�,_M�g����*j_�2 �0�f�Za�������;��������'x�h���I��k(�L:��\8}@|�Q~���'G���z1@J�T>�
jx���Z�I�c��r�R@�F��]�xA�g��'�3�'�koǣ�9�P'�0ma9��a��֮���nׄR2F�N���N��n�4���YzA�w�=�7�&_!� .�m
g����ғP�q�+���&�5��5�ZS~��܄�kvN\�*��Sy�Z��H�:�Zf�H�� � TOo�b��Rc�Y�-p�|�gd%;����!9'B�5�s/Pތ��1�'��n��7�,dL��_���^{�^LH�������T7��}�v��䳟�1�m���3_�;�=���%��߯�G���'�YEv�c�inm��,9U:Gi����;��>d���:��D�d��A��E#��m��|4�#h�*#���!/EM	�:����{��
j�}nE�D� [� 2�s<V"\�yV����i�����"��
{(]�*33u�mFe�MS�+����5[������G7��>�V���cs�]M�r�M՚�X�#�%{ƀe[�)�C?�g�CG����	��tJ�0��ȷPl���1�j��c˻OO� �{�6�m��'�zI����ɤ�%�V�E��6��M��4���x�Z��d���j����e�Ƃ�#Ƅ�-�$/�ST�  �6��"�k!x�E5>�:���g����C
�?��j�� ����.���ݴ��Qu���{W������_0�국�ݕ�H�UdN!�`ÑABO�n�M�pB_?ir��qja�$�Y�!�V�_>ydsK�ٿ}ݭd�)�>7(SEx�@���  D���-�:�-s�$_Q:�wҰ���i��UJk܎~�sWF�AC,ӿx�ٰ=���ͥ�(�Bj�t�`��X�-����-�5(PH�p���-k@�g21]¾�I�ǩY����	-��*\%�/����19�����G�"�bVo����VrV����z�Z! ]�nܷ�	��;�2��E��um�J����e2[��=I���O��5D�6���b��,dIsJ>K`�-=f�}/:
m���erj���{����Kl3��"�ы{����O�}\u;GMʞ��g���s��߂jo��夨_�z��"-5=(��K�M��X��8����o�\Ȓ;��E D#Du���wL�$��r�/�T��b�h�B�y���K��8��������&��SQG*$$f�LQ� �Xf�ri��%V�����9�JY>���P�itC�{6�����z�p#�[S[tד�jqI��ʹm8_@&���$;ӫTG���؀��˝�Ȋ}cX��8�X������{���B?�#|`l�5Ӳ4%s�)G���e���R�h�\�Y��ؿ8��U��u����X2}���C`g�{2$|�j�o4�0]���#Bϗk�FE'�'�X�|ґs��]H�ϴ�e8��l��s���=�7C����#P9g��h�������1��&�F���'�p
Б��	�,z�U=�N �0[�˂ޠ�#�'�n�6���36�xPf/��h���Z�nm�h��wBLB;�gۿ�H�s�x���8���ju���(��F��yc�:�~cV{��������	*�b�_�˪8�t�-�5��8�&QÎ�X�26����i��s��N
>Sd���`��5P�f�7�í��@E\��Q6���-��v�!�
ݥ�K\ލ�Ñ�b*�>AP���s%��X'!0�C����-�0��6�>a�<�	a?���k�2������҆_��,������.~�z�^
ShvQ�"����؉0b �������!,OSkL������o���w����w�۲	[��v�<��{d%�z�v�c|� �����`�"z��@��Ƥ�o�IšmX����[g�e"pC�� x���b�����lЃ���^z���%j�|w!`yƜ������,�i�#�"�u*�x��\gcn
eO��n�Y
��\Q�RS#o��u,���-}�V���	:��� '��-ݠ��k���]CAaբ:���^_��?�h#�#��n=Y�eT�,/"��D\��	r$�<^-~hO4�4*��!��;ʄ{0r��H7P;��>S� �����}נ�5BpW�=���z��VƖN6VT�8_s�'^u�b{�4��ǎ�>�C4h�Rw�+I��)������h� �b�-F��M�����ߎ~�a���R7�v�&�<u�G	Ič�p;&q_rѳ�8F�q~шӄ��B�H-�O"���t��9�%��?m|j��Z�\�R�2���R߸��"$o=����NG��?V<�Rߞݠu*���x��K����0��nz�(�;��$��W�G	�ʷ��,b��1{ ����/��Z2U������w%B|��N^-rދ�K4��\�Q��xDy؃!{�Z׫��_������S����9��~�*����1�z-
s�����b`�L��z�1_����d��m\��(���q;_d$��?���Rr��VE��M*2K]�aiF�'��څ:����(�뾩�+�������yf�:�Rhk׹��3I�V�����b��5�OE@����5Gs�� �X�N��\�_���}�����݅�!;�pI&��&��5�S�r,A�4��1u�7��->��@pX��T!�P�`$�%]M����g��� ����>��7?�t����Ķ��/tȪ��GC�?`b���N���6l<�Go�Wڝ�j��U����*����o���<��e;�z����i_B����F��9�vNs7�Jї�K*�Ћ`?�D ��d3�LA��������ߨ%�����Dz�-ƙ���+�~a��A6�8�#�����|���Ll����|�MX+���,�E�~��ň|��VlUf���k�
S��aӲp����ԡ�������^�b�٧�K��1�)z�
Y֊/�B�͉������;����ʧ_�u��a�YI~[�1����|R��|G�#�M���~�du[�r8��5n���Eض\�h#R�\�ݍQM��!�Qh/V,��%˖��R+��D��0I�i8�jm�!}��%U�ט$yL< l���w�A��"����@훺U��kNM,�yyuڪ���қ�ڞ�g�|m��ޠ��H��W��������t������9X*j�� �ZW�x�j�(�շ�wy�V�b������e�/�IOӰ�Ig+uf��*A [�\@�!$���\k	�߹H\fۖ����*����RJ���d:$RJ=�|}�� �G����&]Kd|�\f�����aa���x(#���ٷP���Q�]�QRe����(� |o�_���	O�H̺�J/��܃��7�C7'�s�#��+@N\����R� u�d�2������F�1��f*)�߰@�kl9�zh���U��iՍI	�~\V�t3�
��F����eVJɌ��x'�'�Z<cw��S��w������P��,HG9�5���0�!�=��\�"%�xx�����-��L�
	��������%z]g�����܋����0+f*eeϪ�
؏�Rr�����05n��𺤛x}�w��!:*��T��.Yt��a�E�w�Ƃ(9m;ۗ4zH����m}I��`�Ix)��KJE�ϐM[�k�R�^�$D�0Ͻ�׊��/������=�#HCO�r%Ľu��Vy�ޙ.��a��
��囘on��\�P���!����0Ć6�:�l���k(s�x2�?x�(�t5���Јu���^�l��8�"ǔ�Ii�#l�a�!(~6��'h����ʹX���&"ت2�o
����&-��U��:�Krdr"R��0��*gʑӂ����z�-�WE�g<��nG�eCq�H�š�<E���Rc���������ͳ��&�t�����Yi_M�0zi"�����&N�|_Ȃ9��j~�n�S�;N�2{�\�Sm���K��"��xF�d����A߱�*5;�&cX5�kN��O���|��]����cz#Z撍V�Eovj��#V�U���e�_����)�[nv�՞bsQ ����G����V��q��	��:�br�3�4�Yg������@~wy[��]�H�n����?�� �2	Qd��}c�("�j#�s��4/p�_��;~PUy��Aq:d�T'6���bwQ�^�PF�A�e*V]R�*�vʑDI?`F;�/��|a�H��Y���]?1@tw�6� ��@[P�D�oN�%^|����e��O&�f;|}�~$"+���_��1�y6��^`<��)��{��PU�zu?ي�k>H�Vx>��O��u�Wӷy2����)Ra�ؼ�
�T��^^�ߚ��o9t3��ʎi� ���Eۋ��k�[l���ڮ��er����˃��r�=�B�w12�r��&B�4�}�	�� ���NZ�������zOU��d1�J^U��D�3��1��� H��\t�q^=�{bؗ�\$�]^��1\����?/3
��������cyqd��$�=����E���y�H�x֭J�	�V/[�=��w6��Q��)�a���|"�rz��?ń)��]�����x�~����40:��O��4�f���o+�T	�ei�G)����}�J��K2�-���-��xm9�M����K�-cvAm�-��d^F���/R����R�}�n�$�k�_1ɡ����dT�L$,_�2�g�	��
6��y2����<U�֜���_�<f�cp7_Ȳ�"qض6�[�)ό�	l��w�e
�� �KX����5`]U<~͂e,ߕ�R�|���ľBp��+�	F����E�K�o'�&w��v,J*q�g����4�Β��q���S�g� U䠧~K�f�N�O�յ=�� �f��X���[����O��([0�h������ �Q4�B|u�9�`��09���wk�����꾡���j�S�%���n�[��91�@���kd2xg�Whg�Q�#�R�Ի�H6�-~{^����0�6I&��^����H�"��GxPчf(��>K����5�s�d'9ڨ�2ŻW[Ҹ$�p��XR�?��^�l���yu��v�����[�h���5.�zm�~휦�1°6y��Ud�>G(�V9���׉Á��B\9S�*	DBt�拢�,{����v�7�yUx�Ε�}u��7�6���1ݹN���#^7`��TJ"U�Gl ��$���.8|֫�ʃ�7�(��������y��]q^��d�D�|�8�]�-��v��'�v׵"z����Y�f�&�T�ڈlaZ��]|Y���Ŭ/�tp8ӟ\[�3�ٛzW �y�ܾZ�'�ݓ�k��i����H��Hܩ�ȏ����{���2�h���������J�;]���eX\_�����.�l��%EXP8�M��O g&�esL0H�4��g�kO��!�l�7�����L!�5��ِHH]�A��'�A�/t"�Ô�1@� W�ݹa�('��ȁ4����J�y�cGůJ`GI!��9)�*��8!^e�"�X����:�jh�U�0������]�P�5 %^2;�aT��%a{@��:1����H�8c���{�9����� D�jw9U!���q�������!�Q�Z�\�i��,��)W�4p*n����1��ʶr#�c��V~:.�O���d��ؤ�+$�_�KZ�(��GBm�'3�����ľ*r�C���nux����V Y0��yXg�!��Uݦ�z�M�d���G�߱�?֞M"��L!n]�����m�ێ���p�5r.���Ù�jw:�se�/|b��u=�aߪe?/��3�]g�J�#���������̄Q�"�
��r#o������s�SX�7��&-f}:{
&�*f*GQ�f���}�{Ė�@{1��>�B"٭�s����"{Q���,�0~j���W���-FJyx�D2�Vw�����"�;V�ـgxq��q���̹�v����Q���|�<����A�y�'%o�o[Ѱp����+`�})*���jn�a4g����Q�'/��W���4�`�7 Yܫ��1��u�T����z3�:�І��Y#n��Q����8W[
��:j`�7o!9 nV��ܠ�n��ZT�/�N38漽F2j^3la);>�.�[�8�4�1з�] ����vΡ���4��� �H��L��[����죈	�g	�"��B��G��~�<�yQ��x! ���nh	�6�u��=:2^�M��5ᐃ�7��r������x�H�o�����(DLvü�aND=�m /o�q�����ʉ��G�We��}6� `���g�S&�7�X+b��Z��ŕ�ձ}*L�F�
�)��!?%�ֳ����Rd��Z� A�db<ީ����1�Ί��Z���cԕӭ��R<^f���t?k�2�Y�17e�����[4�����a�ޑ��q�g�v5Q�K$�+bҢ$�gE㮚��{��5�R�Z���{	�	�D�����(<,J�K����L1�(�W3�<��SX���uoi_�+,����صX|�IZ|Sg�G���1�c�-�'�t�Y��Y����G�����A��z�~�����K��њ������Zt`=�7 '�� w,U����H�z޸�����g��#�Ro,�@��]�Vpv	u9��H.ƺ�H&/���:���j@��oj���{[
8�E\"��������f-�]tZNmB�'��Hm�^M�O�(�`C����=O�?=���@���b)�U���/�m-��_8|�,'>�{���s�=gs�ivJ�s.l�����k��6�����G�)�dl����/������
�*�d�rd2o�{�/�s�X���+������u(;R��I�]g�W���?%��;����6�����!�b��"�q���5g��Sܬ��^�'��2�"��a�Ì�5r7L�(������d2�
���=+�4�2��>�bӦ-��L���l0��z_�p.���_F%-w��T����f��okk��Q�$V�0��-�Zi�]�Di<��YW����ꐐ�t����9"�ί%*?ߗ��"ތҞ���GȨ ӗ�c
v���%�d����'��K��'�3T�Tȹm���ZTB��h,��*|�7��+��o��]b6�U�ըk�x�b�q��˚��V��*Vw#6q�z2��Ge�Y��Ʃ�G��C6�;�k�wM%Ľ�:���5�b3�T�����&��GK��)����j]�\( b1��*��18A�.����Q��7�d�x�Nf��IRӝ�C�{zZ��$�֧��
H�H��Vq��w{���E�le�hO)���l�z\􀤡9}���&f��l���Ѣh��v(�8���@��6�ţꕹ7����rty�:�aÁʳ��dR�������yo�u?sx`�~!�sl��*�"��ieB�3�y��*1�;�ruCݖS]<��-o�j#��D�,ΪwDI�}�c�ur��x$ ���i@B^PWw�DDU���4ӱ�4ǫ���-Ȳ�������Q*[I�g�T�r]��V����s��4�gP�l
KM��0�	����� Y���;�+�+2g�㷻!�k)c�H3Vι�O���p�UK�dY�lYc���%�!���65��6���sy�T�_z1�~)ܻ�$X�{iJ�fbC�Mw�+��/��=�Bя���uo�W}���0x��E���*�|�P�mv
A���	���J�?מּ��W� ����Z�G�0yX����#�.�Nދ��<��0������X2O1gD/u�ڠR:	�����i�'Ȓ�����*�"���Jߺ�/�L�ca�F0�y��?�\�һC�3f��_������ B���jT���5=��]��.&��*�JPqg�32o�}ҝ���+�C<a<hs�5�1�wgc(Z3���:��N}X_kO�e��ND����zg��tp��3�oX�����{������I5i1��^�0�u�PsG�@����/�ɗ��c�̒ �S\���J�S��LRf)��6�2`#ʙn��k�Z��rf2E�l��^G�m4rL6�t	�yP$�ܴ%���ކ�<��*��3���	Y����;��������}ZgnK��C����)�8�Q�r�C!�g=.)꫺.����Ƃ���NtP8�w���L1�ƈ���1Eث���^�w�e��V�Cx]NM�N�Q�i����}��'Y�r�}�t����������*)�u�5����nS�&)������!9-[��#���ő\�=s8D�1�Ұӝ�!F��E�4���=[ �k[`2�r���@+��y�j�Rb�n�`�.P|�;j�#��屰b�/���h�<���<�[�I�(�a����n��Fp���)F+͞x'Ll�zހ��(����(��d��+k�,?��2�^���r%��)\S#H��<DO꼘u��ݧQ�<���J՟O����đ�T����&�!2�������И�"M��-{���. a�M���ផG�*JM����w���G��l��xޢ��ȋr��� ]���$��Dp)��06��g�k��p�&Jg~8��5�q�.Z���V�����d�S�v� ��6�j�Hs� �`��kń^-�$ �ΰu�O6[��R��{]�(��%h�1	d���s>Nz\gAK�[e���<�����2�����2���ȡċ����
7��������rO)�N�������9�s����	��Ӄ��M�榃"�q�%��f�Jj�Q�p�_��E|D���{�?�����R��D��s�_������6v�Տ����@S�"Xt�3�;:���/P��A#�@�OQу@� ����?}y��D��0�"lo&c�|�?ӟ�b �;SKG��gC�,�L�ý�6��e�˸�F�5��7;�!	|s�>j���h�Cي�@B#g[(a#-!�| .f����:�;�ٷ
���%$�0&ߙ{!���S�)O!����=fh��b:B����^oo��V���w���T��i���ͦA�s�"�Ʋ|i�H�����P�(�p�3��M�/����>!�g#�
'��;�y@��C�|�Ս���!�)� Ȇ-.�����|��=��+�u����H���u_A�/	ݤ�Լ��)�'��,C�ʩ�����WRx���H�g<�)��ꇽ�H��k�N?ۍ��]7ha���6��z.̠��Q1���U喝3�/�&/�Sָ���=��9�mn�Y&�l�R��]��!aBIz� ��69�o]�f��.}��v�U��
䤇+߻��r�-2!�x�K�2E7}1�P��x�z��p���30���1mR��+o�K���@�l���Mp�B)�R1JT=A�Z�	6��@LP�fk%J��[K�l�X�7����Z`����{�7nK��s;u[=���Ik�{oR�x����o����2sJ����y��C�Y��횬�ȱ�Ro/��(�:)��}L�R�3���(Ɨ.���3�Gf��_΁���8=���|�'�^��k"v�o@�6���%B�l�א\�N�+���,/<=��Sʠ��j|�D(�pE������}��l���)f�\ 05�����&}��?����2���6/� ��19��Oa�������"���dHZn�h�p�����W��q��P�������Ҟ�J>����Ņn��^Xg�
F�Ւں���<�Wخ�/`I[��$U���۬y(ZT��ڬ�;���מ۫L��y1�A��W~n�{3�1��c�E�gW�������;�䏬��<�)�R�n��N����	C;Ҵ_x��˺-�{�ؠ��Պ����mq� H^�}�}^�̈�Gԁs����~[Aݼz��fp1#��r�ǫHQ1��#x��_knV�1V>"}�96�;� 	��X<���O�u�ljn�(��O8/4�vɞ��o���=������9��(���[Brr~�����"����l��4���+&��;��x��MJ^ �C����%Lڷ���,$M!~��W��%��N�,C��%�T#e%�i-�d�⌝��������<��=x�� ��K!`�E�k��v�(uz���Z���'��P�?���?��8�xR�orS�f��ɓ���l;�+t�T�L2�c��\䙠+�ǒ���߆ƕ�C�/Ԩ*[�!l��]��#��Fn2w�R��ѥW'c�O�鑉��A���hh�#g\��÷`޳��8�,��k��Y:��<�D\�[@��9A�Wږn���'b �v�Qk�uQxO�_�f,u�N�%\���zzT��\�k�`�<�����-J�������V6�A�����׊X'-��oZ[�8��������n<��g�o��sH#Q��մt��g�[OJ�0���i�<2�x��=v�w K~�.���D��Y�U�aS�T]l%)��e0�ڏ�o�@��R�Mg����ǧ�
n{ ��*�����)n�_�B��@������h �i0���7�KlP��]��5r�|�h�) �h��Q����:�R�C.t.'{@�4�[��b7�9୕�G���{�U/u]���u/S������1M��B�ng~P�[p/��g0K�Ir�etE��솕FP��.�|��8���
i;ycp��%9��{1Kg����1��A�&0kd��ᵮ���2 P�9�%g�k�$� �$���~n/9��'�t�f�QS��B�K�HJ�P+�N�<ӏdp��	gL��@��e��7�#R�W�3�*��9���X+��R/Iy��E\ۥs4�}O��#���X�{����D�x{6��9q%G���+]��J4���ᵥz��FF������}G������2�E��t��3UA>C}Ο<j��	C���3�C�S"���d�X����3O���e�fB��q��K����0�T�Ib��9a��a^�R ���3�(!��* U1����+�������&y}!r�CvҚ���w����	��B�T/N�	��yM_���f�<7״�/t�0K�yip�bVr	�X-��ipF:x�9E�j)�G�%ˀ7$){�	�����_9���_�ٸ)�;�ܡ!�Pf���u�/�m��b*%_e�H�L��p|���ym,l���	�!/�]���)�ڒ(�u��-X;�A)ިo:pH�]kVO_Ѽ�����)@uv��r�P5F#���{�5�����	�KM8��}�?*�g�6֠���Q�B��bS�����$�̧��Z�@�#2 �Kp
��@'��@"�B�$�&�U���&('O�~���ߟp =� �-TV�C�|���H%�+7~T��Au����M�qŇB�hm"�`�0C��ғo.~��Iл2����~R;���w�?\ƴ�gЙ�ev�q��CG���汭���P��E��GN7���|�̗ɰ�b�.��/s$�T#�>��3b���?
v�� ps�B��\{��n._����Q��]r�Yn��<L�M��B�o� �y�i�Ĕ�ˉ��]L�9��L8���O���d�Z	cu� ��cg�L|~�ty��̣e��|y��1����ZOؓT�,A;f�XV�(�y�cBT.��>C�����a���	`G`��)Np�3'�l��V���e��fN�b�?YHJ\�%@��(ܬ��!�*�p������v䙮��R[�T8��+��8��2k���DL��ka(�{����4O�(9����L}Ĩt�����dC�A���2���gs,p�kq������,������U�b�u$۷lQJ����Y�É�D��9�f�Hܖ ?Oj�I�ғ��v�c����N˲�T`� ��ј1�1X��U�1n�)��<��V}{zH�Ɗz>-�xtj��H��K��}
>ޚ�`��J��N��F�6�m�zL
F�fhN�O�O��s\&����|<�Ԯ�@tP�m�}�7=�mDFJ�<?�ބ8\+*��ܑ��sU������4G�k��\-�H��)C3G�f�k�Z������}
=��P�s�����8IW�3��J$"<��t��J_�:Hl���都f,��F(�����^����%B*௶a�-Z18o��ҟ5��� 4:��CX]��4Fwub�6vW��0f1��ư�x{ܼ�B�w�����QcJ����k%�N\qzv�bΞ�9a$W/Dڈg�d1��{@��[s��qm�x_�ql����}Y�#^>��F�Z�Ct�1b9k$�r�Y�]b��?E�����Ќ��`�������X^�����H�41h�P�����/V�~���G�&����?'=��4��D+�!^�s���e(RC=�a)��1Ɣ�^1�s�"����n�(�ajsbp%������yMD-�������]-���|�2�e�������s��?�ch
���בi�o�læ����<�ё��v�Dml�4U/Np��A�yS����Z��{g"�#�_=�(n�v�<p��P��F��!7}����_�V��Pm�q��.a�p8L�Uϖ7��Q�2oOL����=��N�RŁ�����T}��&e������4Ϣ���XXGg�R�q��K3���;jT�`n,� k��y0ߢ�f��Fa�~�E�"KM;�����_�����YWBW�,����+)�K/��}'��g깄19��4����4�8K�qa���Ra�+ ��x(� � �:�!�3kS�ZJ �H6��@=m#�n6���	-딦����}����C�|�������4w=�u�����vE��!�ϰ��*[�G'�SL5u�{�d7/�V�,L�@Ϟr>u��l��)�_������C��N� -������d�g-�1����2�6#S`�R��E:�a�]zk��=��煡���O"1����|��$7�T$�s((A�};f$��]�[gM�����m��xY�1[���L��d)oT�c�h�&p���LxO�oq��7k��^"r�����f�~Q�Q��KS"�B!;�B�~W�N��B1�D�����mKՂB�����h�8b�O֊0 �p@����2x�4��p�]2Ѹ�;�e�!:�W��{���{ˈ�M	�bq]�`3:�;I�RDOF���|E7�_��h�!
�(��PI8ǝ���Q6>]�����?�~�sh{p�.��̔�8̓J&�2~��? M�ObE�r���??���=��t��r^��scˎe�k�����[�=~�Ur\��#�±���,�t���c�B38s�^L~h�&�Η"�^��I�:փ�_�mO nBĮ�ǜv�{���@��hpN�cFw��ڠ/G�`��'���gc{e�G(�T� ��!�CM'�j"�P=<1�(z�f�v��+sƞ���#6��M/7�:�������Uq�G��4Ing-���
ц�>��Y�ki) ��K߭V>�xl��>7tp��(M��hlX�fNĆ�!T�i
�LF0T����oO�U�ͮ��=J ����$�7j� o��'i*��d۫}mxF_���۽�Ȟe0����fq��'b�ٛ7]��#�~���{���vW�F-��xE�#��>hg0���w2'c-��Z���|�>���tѓL�3��d��%$��ҹn��r�^�υҟ����;�o^��.19�r�����,%s��v����u�Q�Ʃ�SN�x�׸mA�`ۯ�c�[F�`=�Q��6{xE�ތ+W�Ф.I���w �(͆�Kv���p��d�����z�-K0VeRR���CL���L�w?��V��#/�ḁwX��q�W�'hpu�� y�--�]�,-����������-D�Ƀ�#[�l��?wg��mչ�k�B�`�ڨ�\,���W�aa8P��:e�t�����U�l��� Y<`v��v�O�MI6f���N�vIV�&�G�����V˂8s6z����cQ��6�%iR��D����-��r��3;�O�QCv���۔ɧ j�C�%)����hT�Ui�qm��Fk����<��N�Y':���u5�'-uUt�.V�X�ork�Ɲ\k������ Ī�ŧ�M�5�Y���+\b���~%뢿���n�,}q��=sز30u�l��`�Τ�
�v�z��6H  |��j"��PEndȝ(����ف�P����y�Г��3��LY9ْ�(x��[���+L��|�@G�A��6�MHm��`p�Xz���0�����v��.k�L9��5����j�β���G�c�M9�_\�,f�_�9�3��M���mJ"�������)���>�T��	Q�Sc�+1��o�{���Od��|��6<���/d>������M[��WU��̱�!���h��`�N~d!ό�'�����M�](K~��#3���"곌Ͼ!���T��y-��LdӟZ����2V}���bBR���d�To��_�7�hS�G�O���b��1ygq�r |b��PW����s��������Rkş�"��%��p�~f�YY���u�yΜ�]�N��Od�[��_��9����#*�J��-�,�����H�����FN,��,(��F	ۉ�WrEx��K�b	� ��Qv[��|��H�O�^�e����0�Bh�rg&6��<���qrGI�ųM�w)�
^��ٓT�<.�����������CRUԼy��}�3/YAM�}V2�y���r��qAָ�=}�nȷg+�H�͸:����o�)�!ѻ0j�#��"�r6�r<���)���)�y-c�ȟ�@�a������"��>w���΍�l����=a�Ks�7��~��j����{L'�27E�����*0�*c`�G�����?Õ�}�����ֲ� �"�oO[���
�S��"����4�DU�ʀ
��x�w��\J�k`�F�0�����6��%���~h�k7�ER�(Pk�p��9˸�Xxg�W��C�4 �v��7H�$�b�J.4��b��Ӯ<�����:莒С�6H�Ix窪�����Q�<j+�W|�Ƌ�4h�"�R�#��3¬M��Pc��<�CB�_��xƸ?��P�zj��}5"��Z_�^/�2&�K��13/���.,�r6}���-��y�|�c���h+i�0
_9#f~�2H~5��`���Q�RV�m�A��FG���&�F�{î�u���F�D�/T��~��d� ��ϟ<FFs�Q�@�O.]X��������Y־7���`ə���Iil������f@ �C�lb���L��!��wT�/��Ր�3m�%<(e�$+L��|lZ=Iz�`Mmi>8J.��&�x��]@T�l��\�����V�1�e��=�֟�(k(B8�1:�v2���5�/����������Z��O���ˣ�;JH�i����aGc��<���}���mKVT��FpG84"�?f��#�o
��~����?lEʮ8������9��:uʻ]ґ�����*��(gt��}�tV��*	"�F��# ��#W~��57&adɮ0͗5Ё�V����fˋ�!ߣ��1d����;���֐��ѼD�"�Tu�B��H&��_+S�Sr��-,ԧ��rB��=�<���4���j��L�-��9$��Χ�� �
�>���v�ֺK�GC���oz��D����#�"�T��K��?+J�g��S��,���#���!�`Ӷ����FL��2+� cM�/�N��1d)�v�r�]́\.	���x;��s -z��0Q���2�\H���1\V��;O̎�٫�ï��Ǚ!!
ꔮaA?%R� �1.�42�tD��!l�Yf���[�{e�������L��
�9_Eo��k�ב���=φx_B��O�`c]w��䡏��eS�2`�2�+�WNy3�}DeG�;����I� X��Q����?�2�
�J�S��/ia�2��x��+��Az�nJvh&�edC��Z��z'C�p�+ߐ�d�0�umkAJn���x@71?O�+�&T�4>��޹�5�eՉ]^?h����	(�!n��MP�E���PL`��g�5���ѧʏ����"���E\{�a�),a�=<�_��߫���|�`��8-�*^> G�j"�cJ��|LF̫ze6��g���G6Y�s�Ն�T偁�27)u���*���V#~��$˫U��$E�Ytۙr��d06B��T�p�h�Q�����>tGY�F�I�q��ӝ��⨛t����Y��ӊ����R@�6Ά���ϟh�]�d!O̭i�a̟��l��~t7F�����K"�[��J[�[%f���Đ���yG������G;?|ƀ��~	��xh�U�v����kQ�Xik>���{JlOǴś�\|�Fm��F��HB��RQ��xh�j�J,)cࣾ��2j��Ɂ��訢<�^_m8�y<�,*ǅ����Vf�K�}�;��g�d��Ͳ#��\��t��	[o7"���Ё����0�T�a�FKeD���J�"��|=�U(�Ǟ�]��O�;��5��L`�����E�[;�@��H�n���1���|Q���_T���»�{�(4�P��v�57ZB�U'�{�ޢ���b�|������`L���,�q�ݭY�<[���s�/)�p����w��넌�Z2^-Dz)/c�u�y҈,�0��:+�aV|	V��L����4������"8�e��`�}��a�.�v'Y�3q<�K���17c9#��3��<Q�m����Z=�x�bw�~O^�U�&�ĉ)�׫�&��@�Mv7�A�^L`���^�O(��z�V�{v�uĒEXB���mu�nԕ;
��̼ �X����ȹ�,̪�Y�
a�t%�HC-���G��W�.�J� ���y��3��Ĺ�o�["xc-�s�E���t�0;���h�i�Y!�`��r*��fv�ig���䟶�.�]�����/[����c�Mbd1Ȩ�ve{�&�|��2Or�UR,�n�׊r��ް#���P=@��ʳ�T�F\��
�-���1�u���>��p/��"����go%;uH�L�t�F��g�
��z�x[��c�.�-wMx�s<��Y٬�&�p��3B��qM��/r��"ť���q?�g�J�hG��������ʯ����W7j=����Qw�gO�3UH�/A;wZQ�ދ�e�~/U��n�I��Úʟ��x}��&��T��ݒ��*�QS)�3�]�����;w� ΤsG��n������$�'� 8�s�)��]�ޭk��1˾��0_�"��PC��ȒQ����hd����DY��V��/W��|-�`se���.�+��[	_����F:%[݈@�:�C��z%׊�0>r����W�K�
��@F.�u�]#����P�\�(�P�
���I<崮b0#�G)�^0V��������)�B���JF��s}7N�˷�D�۵����e���ƋqD�T�}���>(.C���/V��]�}��������WD���5��9-���$�P��o��c���/���a�5����(#���,�$2�4՗e�kS Q���=<ʛ_��a�x�~�f��Һ��i�
.�&�QF`����2�$��������G ���~D���24W)K�A&�mL�c��Y�5�kX�;�Sv�
�R�k)��`l0�(sh7���P��7�n��LK"��2qw��7�����b�G��hm>j����u�v���h���@��b����_v`����N`��C��xE}���lx:q˃Ei��B�i��-�u>�8�gkez&^���<P]!L�LZ��s��J*9P�nGvd���6Y�����{�{�'�	5UZA:MJ�%r�A��:+:��N�{�[_|j�3�a�3�)44A\�_��g���DH>�"����5���%�5*$�5�́˶o�c�}�d�e�b�����j����3��G�_�����2a����w�>6�꓇�1/{�-��N��Q�<e$�f��b��c"�k�t��<�����P��"�s�p5�	���Gaz[չ���y��t�u�[�LE���Џ�	�a��_'|�"��Y<�-�Ff�����
�Ր�J��놞m#Rv�	�K@���A��{�!d�6Ф�������N��R�oj{<�\����1F=e�@iq�_���J �)�����z��?��f�7L�MD��N�������J���e �A�^W�{|	�\B��ݢ��E�Hd`���!8�y���H9@�$�j����0�u��?��ӡ�J��j����.��I�����j������i��@�ϼ�{9sc����pף�����8'a;�dg"W��ԃ���m÷o���?�1]��V�9��E�3�_q�Έm��=���]"�y�R� A���[S�zҰO�J��ˈ��c��������^�S]��cnk����<�No�y!�p�'������>��`�E�\��6Kpk���S�&�ȋ�����w����1�N���Y�􄻸�s��v�v��w4]�ǋeF����PTe�D5�!ˍʱ\��ǁ���=m���B;sU���x��ϟ""�g�����O|b� ��W`׺��ߌ��Ԯ]4�A̰�2��h혤�;�0d�jc&��*����φ$ �������]Q�3�����|
�vs;U��T���V7�����lI¾	�Բ߃��΋��G��ϷP��%;|�״�P`ƞ"!Wx?_� �@�#0s]�����A<v�_��Gk����N�����lQX5���Ӕ�ٍ*uW��,���Q�cZx!�LT_�r�4I�O�[㔍�?;,p\�8�Z��3L���~A��u���+{zg���>%)�_�ft�UI^Z+{d��R\�K�LO��R3�tX���3�Q���2͑�1#@���ג�S�E,��@,���J�qb��|��y��)\.IGOn��G[�����Q�MXNh���3�fS�F5݅1jS��XQc_�js��x!D���^i��%��%)(R �	/z�j�����E��~�:<_����A�[�@�ܵ�P;�ߥ(�s�`�)�5��y֠����7S��	j1��g��/k��jDq���S/� ���v����o�����Ar%F�Ǆm*�J{c�	��ĺ�S�G�0�~L��S�9��Ѧ�$��Ta���:�,�v�[�%'���	�L�ޟ�f�{�}��\�]y}*�f3\}U/}c��"3?�Y�o�r9ٲ2�)R�,�9��h9p�����:�0��Z	�h�4D1^�M՟FxL��'�?]�A�����8F�\2g�O�~4cD54�[�2�[�_��$�G4�E	�=����0��X����E��� Cv��*;�S{�4�)h�Z�����w ���e��i� `n�
�2!�P:�kO�r��J8h�_��*֛aR�%,z9U�bj�%"�+]��� \ׄ���N�䗾.z�l��񳲖��M�v��N�����1s§|��mA��5L�gkзF�M�Z�I�}�PFI9��ey�D��".*�	��(|w��X���V[t, �*��]әm�4wtl�Q8'�@X���2Z�AMx4~W?���L���ƙ�w2h�����فօ�B	��S�􆿄�DMW��,e	��k��▝)�������V���py�pNl̋h�mv�U��q�IW��u'�3��Bʢ��J��^�'1�����u{��>�,~�䌚T��K�h��)쟯 �iQe�k=ʏ���QRR����c��������	$�[�����^z'�����y��V�#��i�i�/��{N��)��E�)1�������'A!��nڟ�n���o~w�Cf �����3qbD�+�ZMd8�ncb�� tc3�]WB�*Z�YQ��LGl@�8K=�k�C��Ξ�W�Wu@J�y�>BB��6��)|	S��x�dv�Ne�GJ>T!��"���G��p:��jQȎ���_��ֽ�8>fv�s��v�XbX�q��h-.��b f��f�Lf�98�5�5'�����1!��ı�}w8���]Y$���d}<�SADn�)�ܶ,��S9�4s¬����<��725�֍D��<k����n�m��  WƑ��ݛ����J��]�7n.���gwiZ_��{&��.11��,����8v�������5�%���fyU	]��T�i}�~���cS�$��´���g�E�Az���*��Jt�K9&� �oDL��P�������;�ژa5_Fu���J���S��nb�N��7��XE~Q����J��c�d�G���:�h�����@>@붰����Q'1��R�nÙ%_)&��3r�3G����Y���e ,�Yz0M�rв(�7x�7�dl��D�)0[��):40[Z[�RN��A��]?p�D^W+��W��U�'/�y"�����F�I���s�_�į�K�d��	K���#���r�y1E.�͆���_,�kK�] X\�k��i�9�c CȦA%��8%�>"��^�}�D�(��!�m����Y�Ue�Q�b���4ɔzMw�<6fΛH��<������/�~�Y�����8�=+!��+��gV�1N�c�:X�A=d�m�t��1�+����`3��(���B�_G2(���W��}3�0a~>���ލ�q� �c=�i�8~
����wH����z1���e4�C�^�������c�G��^�G�WPr�s�F���3q�Ba��a�_p<�Y��]w(�r͑���[B3���Ps� �6���k���-�U�L� ��)u�DS�;�/�'��|���8��Fh7�+Z_3H������5�*{�8�	�o��Wf|�8"��N{��>e������������+�
��b���Q��$ ��)3�& � [����س��1��U�@��%���d��0�p8�j8]t@1�ࣻ��i�N���MW�<M�*���>��ŝWED��d� Xy�!e2���&]\(o�-_?Wؖ�&�oey^��l3�V��ʪ�4��&Ѳv`���E �_��%�aFq��'��kP��cO�Y' � ��zXSnG���������W���~Qcī y�����Yw2�~�'��X�N���5�1�P�\�A��0��V�Po����Y1�%���^��g��"�\q���7i4����z
r�^ƪU��A%���v�k2B}b1���� J^�Ə�ʑw��v[\b���]���8���
��Qh\��Dɶ���?�7�&������	�s�^9�\�"2z��27�Y����5�ث6r�c���K_
Y���1i���3�Lz���&#�O�F��$b������t�xg��U���
ܠ��X�M��_1Hz0��@$�
 j��p.QB�J�Z�\�D2�&�/;e]þ�>@/,��a���ߝsӃWڊc���P ߜ�1�<���-)��:�.�R�C��]��N�E� �ೄ0���;V�Q3��SˋǓJ>w�k�d��}p�V������@�N��/Ŵ.&�l�o@�] 5K��?9���5}���G �Ća�e�/���뚅WR��Jv��\�<�S&�&�D�E�fM��r��]��*��3џ;�ƆY��������W�E�������AH�&�ɰ=>t�]�κ̞-8xq�̨��f��Q���>P�#�o����".H��$�ӹ�4=	��s�*o����. l�~q�Ku���C��di���j�=�����8�U���J�����b�F���:����5�6]�iN*�x���ni16�JQ�����1��ݍ����"���){�y�� ��N�xs�����]L2�Hϟ�"��
"�fX-�֧x
<槐P��H�v2q�Bt<�Q�e"���^tH#�2{ �Y��-9�e�{[Q52�s��H�ѵ*�W�����h[YV���bvQ��q�;�q�j��B\�k�����^I�������̎�k�ӎ�*� i��&��vTf��ʘ��y�{HD}��A��8U��Q`fR���_����m�+�3.��`*8&��Þ��8�RE�uٟ�3��<�7�	�u����;��L����B�5�>����
����h��5A%�CP#+��s�x���$��,��]��}��<"\)��Z�~�h��W] ����>H-���@�s��
�Y�m[�G��{��E}Å�"��5К%)u��z���~)G=���>	��}b� ��v(�.�7��kt�*����a������Mr��ý0hC�k ����52d�R�ޤ��lG��>p��w��t1g)W"�p/<�ݑ
*���xH� %�l6����srH�Z-�ˆ�b��C�>��3��Np)���i���\r��|����|T�ԩ����ט�Gr޲=P��a�0��9:[]��^�~lP�zˣ�^�,��/܀`��E��D�s%�Tg{�ħ�i��U���:�����0�uC�z�T�<P;6k-.oTZN�gx=JM*�=�ų\�eݍ���W7L2>ǝ�^RU[��'`�;������1���P���-��R�*'�7�q����R����m#�?�Σ����d�돰��ݕ���C�`FFQ	.Ĳ�Q�'K҆Lɱm�� *2��:��hv���d�ص�΀��~/L|�sV�,8���	�����&�<0T��u*���L�3��!V䍂Ɨ��%ʺ�m���x�
�����|�!�dٿr�u���n���MН�D`��
��Aa}3�M�>�aجޭ���p��*8]$Xs���3s]uI�R,Ջ�O�V�A�>��I���Q������P�z5�%����es;i'}��A�'���|/�Fa貿��ѯH#CSt7��6	f$cE}����%,	íqi��V��/C�����mA�AB��L
P��$5�W�(��a����Z�a��}:ݑ����x�@q��r}�`�U�+��t��H#ن3ɢ�8��=��ۼ��m	i�����$8f'�w�ǂ;�sk��;�DεŚؕ%׾0g�Fo Ea�0曾���>�gai��<���
#����>�^��z7�J��/����!�k�Uy^SZ-w'�ĵ�.]����I���ua������x���&��u�)V孁�~x�X��D�a�͡�/�w��꩖�߄
#>۟��}:�e�ѕ�ju�p�.��T�b����4�v�0��ϫ�䝋]��I�ߓ�k�Q���C�A���3�?q>p�fTtsy E����Iu�$�R�����b~��%ۺM�:lb�uS�3�.��¤n��K�;IC^�C:|=*t=���9?�1��rؕ>��������#�2dɼ�W�?)M���/6�s�;U,Cp�4�®ޟ������_Ȗ�����YE�\�K�񕛂+��5��%��ܸ��&��i+��k����Fv@P�Dt�3����
I�ƍf9�#䄄�Tʿ$�ɨ�+��2���V�������7p3�V����yE2��"����]m��Mgy��i �%���&��dq���\����|��DH����+�^�9���J����� �e�u6��I���1p���w�7��09mt>�\��As���1�!�S�N)Jٚ�+�e����E�@I3�R�NEl
6��s��Q(|�����}�����Ã0�F\aG�p���:����|"(�(J�u|6)�8\̐�L1g�{y���<�ȯ��؅�|����^��-�ne@��ߧp�B�\־+�t���6y��)�8�n�ci^6.n�l!X%�mR�RǗ��bו��#y��s`��vƯ��]Z�$eIWbeF��ּU7�����rl����~gI�7@��..������:xRbڟ\>�	�O7�J�+^L��D^������6E�k�L�����1�z/�u<��+1$��5lcZ�4�ކ�x��;<�O�F��YaB�YuQ�2���6dj�n�l0��-���[b��`���|M�\'aeZ��O�gi��s��]��ex��'f�?C����&-���w�,�=K�1�Lٸ/�ҡob�Wzoѕ�=�k�9Q�xql�>0��7
֓�~Rrk�6I��c��*T!�1��Z��j�m�Б�l%	���-�&�f�^ʘ�-�l�n��y5���y<Y�9�6� E7�hd�� ��n)|�=�b�w�Cm'2F,L�Eꗼ�>m�jT�����+p�J�ϨI$��5E�e�}����-�)�h�,6?�qP��;a���H؞< tZS�ߎ�ei8���A�[��nZ{�|J)N8�4��<��E�J#��-��RP�u���V�����׸��0���N1�R�vkFb�u�z��"�禛@����;�f��5d��ҵ��|����r���(;M������=dm������f� x�&=��)��'���0m`ɉ�g��)Yh4?
��D'_ˊzN��)VH�s�"_0�6cR��j���Ro`�;�$M�u��c>cÏ��q}Q9�����P̀��Jn���qF��2�UFߒ~�ӝϥ��;>
��*yx��8GŨ����Ƞ�A�~̂�M��v�'�)a#����n � �?E��_�b!<�nr�
!��Ͻ���ш���Ϙ���j��6�T�޲�p����
�i�����}y��Rԅ��l��u�J�:�|+0�ܔ�Zܱ~[Hj��-lT����k:���n ����� Ѓ�"
ti�hV
��ˉ��5L��m��wLϾ7�+<�~޺o�%8.v �e�W��|K+!�<���i6$�c���ڥ�0��aɟ�����������*pۚ*��y���(��/�An�%��t�
�Q�fo!*�Hb58Ѭ�/כ�����#�@rC�6�Z��ܤ�Ǡɛ$�rP) @j�}�P�Ȍj�� ���Խ
��������Ƌ�{K�X�U�7㵔��|���#`������K����%�@��U|���u� �_�hl>2���{�gK}W\yU�vm�����2�r��ʕ��-�Ͷ��*����VsʦsX��[M�X��;&�pِr>DQՀd��
��Y����V�]�"E<!�S�} �F�j���K��䖪\5�y&數��T�kѰR(JR�V�����L|���[+91E� �j,��	L`��?�T�m?�ŏ�RR�%`��B*���fߎuZ�bF���d���h4��?�z�&������2�TxN���j�a�@	�]� d$��}�)�G�9��/̂�p��k���1�5-��ek3W��蟰%��{���?������� ��#�̴B���,��jî��IG�W�g��wB�9�_�oR�͐���E=�۴��6�D�U�Kö�N37b�޾���!��e+������jyH��e0������s�^\� �E��.���v�.�����ZZL+NЙjp��K/����<���D5�Zy�{h�R��p��<�"����T�j���Hq�Qk|ҟ�&�;6R7C�}7�-,w8�e����(�~�h?�u*��n�v}:}a'7�-����^�]��K���Z�:��!�rm� �]0�\6�$��o��a|���ѻ�}�~M0CJz-x(��]���h(2�5*�PgA��kP`*�c
�0�$�c߸�ܶP�m���hz�ʠNB�NQ8�Hb����ؚ���S R��� $f�`���
S�Ƙr.��So�:VN����:	_��]�d;/3s�Ю6��	��n,^���|�db��T�B�صG��p]΍Y�b���-�B���[IA7I���k�q�ab2	�uMK|�����V�~�݄��.���C0��cI�jk~�1�g��7�zc� ���|	���o�k̟&'�O��9�=��x,ފIK�.Ĝ�OJ�����j����D�l@�Ngf�6�ŀo����UFP��+�8�����k�pl�Qp�{֥~����w�}����Uro��'{��IO49������Kcd5+Z���۹��zZP�a�E� ��E����/5X��4I�ƍ��kigy(�SD�+���Ā9�g����*���8(�VB��.;x�Lǯ��~=�L���Gh�c"�ٽ .��w�u�����&��"V��2���,*�����d
�~��[W���M�@G����̐IY���0�b����֙�K��е�:�fU�?���uL�Bs��eWn���.��C�&f1r-4hE)���I�<��QH_HQ��$��Q�)����c�m:�������u����OŒ6� i)��c��c,fY�t��B�eN>�8�|����V�m�y���#��[/2� ��qpq�Q��S+��/��	�Б7,St B�?A�q\3iN��O}]èR�f��t�d%����3��*˕eX�����Ԑ���K:t+g��Ce��ZJ��ԿE�FZ�
5*�P�NT�e�����[M�1c��<65�v��ȴ�:��XA��O��	=�$��D�J'9$�7f$~m�9��UT�L�����$�V�0�w�� o͖�b�Ԋz�lN+�F��'��q�}�>I8Ry���j<{\9����^		n�o�ufA<^Y?��{��8��h���\��_J|,&f�����&���&?S�r�5�Ԕ,��,O[��o>�/�\����*|�v]�\{��Y���}�Q2�I	k��[�ڐ{�
�٘R�i��oc�r�N��~���`wݤu��1�Ԟm��@���Do)Esu\f�vʔ,c�����n׷4�iX�jK���U��+'��� r��KȲb�K�];>g��
�n�I;�J��$$fݩ.�4�?�N7�Ԩ���D�<H�曤��bQ~>!d&L
}eq�:͋R��Z^3�7�q!+
���Ap�fCm�� �0
�DO��BX�P�8�|���~5j~>� b눩T�D��8����*������C8t�� �x�O7>ƅ�a!�����k�`_��,�4�E,YTD0V�4�����#^��?���0�UT|!MB�/�z����|��K�z��wc�}>5/p�`���$y�"����)��*#���:���_2Y����k���Zbi8����ksKiV�