��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a���?�;��ȎɌ�K�-B���b��Ƚ�/'��{��> ��	^FV�X�;^iQ;
x��}3�X�R��/�b#�x��*�"xH���M���'NX�䕇�,�{��m�D�\�%ߥ�$�Lo�:htuR��$E$�! ,��gm�:6F��1%JC�� ���uwJH�I�"w�e����o}H�Qʿ@'�1��k�l�ÊF
�G1����4�c̓�u�c�E	�Ԙp�r�|�a���w�7j�n
�n	�	������b�Q�����x����!09�\.K�ݩ��Ǳ�.U��9{��b@ʠ��A{Y�� *�usMZM��0q��:mޢAЯ�)�+��I���5�=6���Y�S�e|Zǧ/��:�!&W�wg�� Y�}�$�[�	�b�~��Q�zZ�pOJ�B��ݳ�(r��PHj��@�y����-X	�v70��Y&�8e���ݐ�`�'�[, �������,��K@D/��8!�����@j�6��+ţ��yp�����qh���+�J^�J*j�X���d+�j�'F��l�5[z�!����dnAe�����%QCS �L40k��據 ���$�9aȣ��nw���yY��oܬI6�*��a�����8-��mqo�x�)�5)��Z}C�h�D.]�Ptr+w7���ь�R�$����G�׷�Lpe:�kS�h¤)� VR�(�O��)l1�b���⍙#=)q��Wz��˿���)���d��
�h�S(T����;/?���G��/ɗ��+nW����3��	�g,2o��Q�}m<ڡ1��nz�ǻ1�ڴy��D���Ծ�"�(�f�VY�s ڍ�yY�pՇ��d4�r��\2P�b!hk��4�N� �ڏcQy�]�M����� ��Emy�lE��>,作a��b�Ch��Ō8uϹ�#������2�L_jU\	�/n!B◻Mt��%��K� �8兂++�d6��U��i�Q`",Y|r���U���V����l�_׭�3�f~�l�_U�x��0�F���%�����?��v�G�,	:��!ܧ�Y�a�}2�168�;05���΢��8�7y�e!����s����*���T�� y�\��<��.���4�1O��z�6�m��N�<�W�����зvx"�z�2GVTs0�T�6I��{�6c�lXN�A����w�a�\Gd+�)yH��R��ee?�tW����yAC�?6�ek�4��~��D'��X5�Mӎ7b2b�e�Jؙ�;��>_����6�߇�%1`G��{&���L:C�&����jQ�8an�`���'�!;`iR�?�1AAp!hf��'!颜����ˢ�n�nu���)��挿Bh�]-�?假����}������`L��|�A�Gܜ�o�e$̏�#P�ֵ�� �m��o/*�5Wp/Y�ǴSϬ�s�/{tGf��V��sH7�<l�/A�Қ����Gg�I�w�it��)���e4�_�h�|��E&�b���dkd��A���Rա�p�	fLxsN��#���;��ŻZ���:����~��Ue��?e���px9"��ӏ��H�������0�y�w�w��������`˳�V�l���\$���]�L��]�y(afDʴ�P�Q饧�Ϥ��E:��0LL�,����� �)A_{3w Y7��#��vК\��4>Vg�>�>�7ks�|�	�D�:�5Q��&<zl'N`�d�R�c��4�3�H��A$p�jR��s`s.o��9�MІ�ԑ+_W�@�2�h��n�p��$��ڛ�#;��N�A����a:M�YR
f�NFjEk�u�$� ��e����;����X�s�y�q��A;�̻BnS�߃��m�<�3n���3���FZ] ��>�����T\��1��Pݜ�	UFJ�WD�}c�y�s��$�b��WUR��ׇ��(�������I���D�>��5��Y�r�>�{L=M�ULwA����f�Us�KN"�A�@��'����>�N�xZ����	�W��]�9����
y��o���:��������v�	���xXjr34� a�C�͑��� *�!2��H����:�ӊ��v=����qQ����#�p�S����\!�C�@ˎ.��B��{d�*Ҭ�ގ� �h��_(���[����E���Q���ȎDk?]	D�9��=�_�Iz�E�!^�Uj&�[@N��A�3�Y�L[�U� w�y�٘������`���.�32�>Iv�f8�U���C�����?�+,Dd�"[<;��=J��o1_�:��]ɛw53�"MM�M�'�c˯q�/���ƼP�&����#f,qWw�fg���g����&���E|7�+��,	�L1��R�j�"x�ߔ��7x�uhj��V�7�̶�fy�&�x%ǭ��P���/�p	�h��d�%Nhe�s�E&��N�E����z��X	���gY�����@��"�hs��\�b���r,t��,Bà��T���;,�Ufp$ǡ܈�6�{���ԏ���Ʌ��V��|��u�mr4��3���Ep���@ѮH�]�#���̯l*��m���f8,�GB��dǦ�y�z#`���'*1U�w�^�ƭ+�F��t3����[qٿ0lz4�B�x7�iTS4-_m_~����xթ~��׺�k"f��6����C�(#s�R�H�ӹ�1��T��ټ[�t`��#�B�����5�	P��+_FU�Ρ��o��/���������-��p~m�/�����ͤ�����x����v"P�d�}^%A���`���z�i5�!g��HǻW�
�s�}�YA�7Tٲ��\w����N&��EhSв�nq}{N�֠oN!�QH%t���8����Z�A?z~�0�k4F�O-/.ׄ�8�
��,(�0�;eL�+,�'T��R�{-���q�]#��Y����\�w�gzl;�yN��PH��f���	ȏ�¥R�,�#������.�.��\�>h!�����M�� ���mS��];���}`��t��QvOoa>��9��!�~��-dv���b0��#A`W���#<ŠZ�Y��_�>���s��ub�rw��Q,�5�9a|