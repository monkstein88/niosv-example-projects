��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a�����{������#��j��{��	?+�g��-��"XSʌb������;�b���/��.v���9�Cr� x�B ��q���mL)�-�"6|��hHwg��	��j������猽?�����?�__��n$ԗ�����NÀ�-
�R�6�d��v�����t;��df�!�+#G��Բ��87E�1�R�x��)O�+�w�v\�A�B�i�y_7V)�5`�@uș����J��E��9zuS�H5U���	�#�%����BV��_!&��jf!���ٮ�rSe���&i��A-xr���9�}�οl�bpP�	��rI��ɶ����FO���V����� ��B��F'ge/��uy��
/�+�냛�gn��+��������_�Ńq�\��(	�Lר�Y��T3%M�������@�҃J�����c����0��A!����d������055���)
h�� �4/����8�M��JT<.�nɷ��:�m�>k�B�s�(
zʣ.R6�$c�/^Y�����������:��� �㖱�,*/`f"�=;���Y��W:*�=$��m �T.���Dأr�����GEi�j��t�ꬃ�/�:%��KХyrL[�k�~�^�����`i�0I�¯���Mu�ﮍ�+Q`�\�F�"f?,�kT��ľ�I�m�}-��؍�#��Z�:Sܞ�C�̨��bЗA�B�b�iye`�jH�n�B�0}�_�!ȕ�~d�����7- rI���m��Z��g�����;5"�Z����̓i ��3����eD�j�����+�ni�լJ%g�QT�8d���`�Mz+�?�AI��������X�I������d���<�G�:/A�� ��{ �P��e%���ߐ���ٝ�  ��9�h�k ;�u#t��ù�*��/^�k�kት9�2.$�A�[�u�P'�8�Tfˬ�`z��2)�>*;� Z���a�!E�X�s��b�d�Ę��寘�qt�Y���� m���jLs��ٖ�A�zk��n�>���w1w�LPh�
ֽD�
��
'������̙�Pyp�q�H���hB>��[��7Ud	1�wރ3�uQ�1�WR}����ul��;�S�G�Ю�nƗ����щ�к�_��d{��=C�d�!����pz%]S�%��	�"4�݈�n���B�U��6�Z��_������UD��%ɍ`U��w�}P�3���?X��i��u�[�??�&'�h-Έ�56Z��u$v����&ד�F�x~q���c�u�
!zu� zY�g�W�+��ǹ��!�-��o��3����fZx� �L��"`�a���I�!��H��}��P��Hf��$��*���������dZ��u���f�I�J�x�����d畦h��di^?N����i����+	P}2{aP�.ņ�f��l�2�Y���ʝ%��v��;!�^%�X�o�X�<#��� ����OzV�mf�Cy�����k@���-?;�KJ�餪���O���x	�hyZ*6܆]w
kDx[�2�;L�%n�˽Fٵ
���-��ڶ�5�~�<�9��}�ե	��9O{/����p\���'�E�k?D��b5��.S怒��a˕w�{?�UYU	:z�*{�vqۿ���J�wu���y�:宻�(J2/��Gu�hY��ϭkR������4�x7J���;j�unq�C+�J���Ί�4pΞ�M*���E���+�E����ϱ"���P�����}�
JYV���y��$:�����&��G�Mm<ׅ��@�ɯ6-� r�`sZW��f��bM���(���Mp�{࿔ŝ�t���;��Ѹf��&�Uʯ`^���4���LI���n8�u5��[�=xj3XJ�#vȈ�%X��\�|��t����DMeD���p�?�h�ftlt��ـqN٩�8P�T��.�0�X��Ʉ0� :#�^����s�	�AA������%�v�" �(,o]wv�I/���$Uç��p�e��w1�:�)�x��K8���"������)4�Ի���}�s%B]�Z�s��&���>�~�;_��w����?N���br��J��R����ߚ��v�q������*�7't${�MS�8�K9E=9�M�u��v�|Z�,���B�� y���pq�#�e%�٥��+���%��K���iƥ��Ö�Z�ΘB6�N��\�L��;TqX���?[$![M�aV��TYzK��9�z�;v~qh�i��߅-�Q��#n�$ S�y\���^���<�V;CC���u|�e �=6%�'��0Ъ`����_��0�C��_�q���s��mKڬ/F�����9�K.Ȑ	(����F�[���)����n� ����n�Hc��l��� �V�¿凂@?7�h?�CIS�#}�c�⫃�Q�|� (�6�̷���qN�zP�K��s?������Gwk��j���[���_��8��vw���&�\"=I�6�/˜�4z�!���l`�Vi�\{��N2TujX����eI�|3sY��<��/��7�q[�q�Q�#����DlË�m�J�LI�\/=om��`� �6�i���=�T�N�2gR�JՌ�s1����d�Y�a�
OT�a�@�G�W��b3��\ƺ.�l���4~�f���p���Q0��C���u���8u��D��Q����-�x�P��EۂJ����})���tڇ��\Ę9��ͯ�-e�P��{L��{��2�Péu{D�wڇ�<
�ՊV�V��M��=˕#�*�j5���pH��d�C��jl�a{c����42���*�ܳ(�k�@g>Ǣ��V��u#g�E��m
edHH�S����Ȩp��zXF�sP+��ov�r֐���z�/�Bv��ymؒE�;hq��s�7"504���:n�$��n{�|L��z���H�-�3�RC��]7�Ġ�(�;5���;�#��|��ZHP㬤�2���d,��Qk�{؛v�VWO�89[Т�:}�@��$����n&?6�k�Pva�ulM#�3���p*m�̝���qY0>�=x�R/%��ٖ�`��`��i�iZ�:]���su~3����#:�E�d����Y��;ٍ5�/��3O��MI�䱃x� N��c!|I��ŋ)��E.O��|[��h��BWNn,�{������_��'��3������T@�nQ=Bo�C�y�eL�ehi���/��/������@GV}u+�\� �,3�Ȅ����x�Y;�)e�Cf�/�Q��=�������j�#���=MV��e�^��Z�"{$�i�s5\ͽ����ƺ	���<J��j�N�pC��6+�6r��<������Y�S��C�4�c�i�*�9��[��{��?po%ؽ�x������K��=��Bz�dL����Ҷ+���t'�(9 FV��y� ��l��V���hC�Q��J��G=�̷�X���u��͚�V�9[`��)��Q7z����4&�Tx�U��O��-
7�25�1�+�����z� O&��T��O	T����6�%���4-C��~߄(��㼊��u��@�,�8
>�7*ڲp��D�-E���D��Ф}��2�y�*-)]~���R��/�D��m����s�DK�p�e[���ذ`?"������
�ί��c_Kߟ�f����5В~��S'F�I�Gt/[�z+귾��×%���SG��k��eƊ�v�~��;8��+�NC'M���;r�7��| �k[�9���{g
���*��_(��A�E���V���� �,3���*��(_j�;���2A6j���~Ou��im��F���t�݁+Q=��3���*�ȣK��Gh��-Y[�0AJ�{>1��&�2W4��܄ǀ���ED/��͉�eL+G��7�Tr�W�-�{��8�d���o>n8"p|~È�0����c5s���m��X�Ȉ�/��)���հQq&G\��趌�/݉읯zI���\ P�=���B*h��-
o��az	�  g��+�R ��B:Kg��ʁ��f[q �)ǚzPa�NB8G��G�� C^]�zN�i���,��i�*����|॔�D���`��B��<�-KEj��$���! d|��vqΤ��	�;��(:��O�^���O�B��
��ߛc;N�T@���/�4p_��7���Z��P���sy'qp���Mq����O��|�˰���5A�]$6LF�SI��&�tlt���1� �5-~!p�V�`����A�s�8��^F�cN����������=���!]?p܎#0����`�L~��O������R�j�:��w/��0�ApO��!�9VIՇ�m�Bc���̤�Sc����O{�R�HE.w�k܅�L�D��@�)�э��}� ��>�c�2d9'*"�vcb��ݻ3����/j����׋x���_ȣ�`A9�}G�Es�Y���jj��
#����6�Nk���I�Y�t��qޗ/����?�����噊�@zi�/�\<}Dc�|�_��x��j���N��E��=X�7;�����cQV⌗�����X\���<!�6ณE�������l�2��jo|�i�0�j��ᯐ��\�qJ����V9��c&����F%�S�]��@�9�:�o?�%alB�+��{ַPJ/@���=�㚎fCmXl�d%l��I��`w%rZ��mL%]xŷ�����]4I� ĢP�F��ͣ�0=�G#��7)�!zٕ5�7�MG*8��?=�J#l(�G�i�X���e5��o��ӵ���5�W��A�Bјy�"��%ܻ���h��⏇͆"���_��罵���ٶ8�Z���6����(��t���D��*�-���P�BSڟw�T�o%�Jn�KK�r։�����5�q�Nj�N-(8�g=��F���(o��n��.czѧ	��5N�&7�k.v�e2��di�qch�_4Lm!����rt���r4�|ꅻ���e��Qφ'e��lXJ�ft�P�N�G=��l��k$�X�N�����U������9!�Y=��NF���[E���_ܞ�h�~~�H�+]3$LCm��hżJ�����a���/#�9�RYan��چ��dlm<��xٓ�5�ff�Ei�Q��U��N❭B�$�����!�Zsi��������\a�>F�)&�f.*��2j!V@��l'GbY���|���r���q#e�QU}�B0e|���%g�^q���G(���d��
E�1퓰�թ(�^^����2&Mښ�K�X2�T�-��yM�	$L�3�3Xܲ�,�������J�Wg����O���>���8������v��2(�1����ӱ{��/�"�U%H>jy�-y�7��K�d8�R��oW��T>1'����7���֧�,w��'@����2yo߀9!o�w�T��ǒ-��& R1��:�[{����f�M��`��	-iw���u.����.��� �Gb1�#@��A`��OXr�hy�LY�����L���B��n�g�@��\�����]�#ƃ hH������^�q�a�)�qY�>���b]���R8Ʌ2ĩ�	�:��;?}s�8���ѳ��#���" �U��̱�������b�J>�8�M�ӊ�����D7��%�?��P=j2�آD�1�M8�k�z����3*�w��˟?]:�)1��f��o����ք�Hj��$��������#E���d��'��u̷�H�&� ?{	ŦS��O\�����
�ׯz1���Ҭ��x�ѥ�sGRq&:�B�g����T9�/B�A>e�3~���ʑ� �ӓ1ڲ��n
�n�3�E�`�"i_u�����26;��_Wy���wv�.�ه�p�u�B?(��WR}T!���Yn2��E�Ms�_�=��/���S`�DF�������m2���ƛ�l�!k�� K�յ�����͕����*��aS��ZJ�@Z�����������I��Y��u!���lհ$��6������6�73[�(tj�;�,
_�5.��T�FFt�+"�l�4��K�8!z�����T���|�ϐ|��0���JÕ��/�� ����桦~�-v��y�J1���/�#����3����PX��V�{�{�׽d\L�����y!�h-��DL��9Y�e�l �_��K�u�i�L%�ش^��˳s�e�c{T+xM�$cS�c�;zkUV/j�z_ �����V��H-� ��r���ޒt[�T�B�&�S�D/�\f�#����xh�}_5�Ϥ�pgIc�"!u'���k#�$�Z�^W}���/rXv�OP�!f����%-g�A��ֈ�D��v�� �����b����H�F�����A?�������.����r�G�L�P2b�_CV�D�;�;�;]�7rͅ6r��0"O~^>�d�������0Y�.`J���:��,� ���ұ*�S�/s��X5GwB��:2�g���+i�Icc(�'3[5��b��&ԑ��w�^�B����\a\a�f9�?D��[j\���f�
ZSGu\*�=U�؊�:���K@��J�W�&�˵:M\U%m���у�A\|�Jx�-4��>�́�EV��I_RZ��]c�=��8����Ye
VЌ-<dӾ��/ �1�\v1�G��R����#>��
��@>ˎ��E4!v��Z��9��y�]^�F��6�h��>-�~m�_�SWє�4_���xk~��E��\1���R�)�	9S��I�lpσ�i�IC���[o� 0����:�϶�����5,�|2�*M⭟�e�5�̙�cu�B��n�W����-���� �C6~��d�Fk���x��bw;w�����$�M���C���7�#��I�Пa���Dg�¥�xH+!�Y�</abR]V8شT��'A��Y�!�e�)Y���3<TC@�l�w��7~j�D8�,�h ��Zw w|D||�.iO���p4�Q���� ��c�אk���I�#\�<���VM�&X��)@�Ax���e�@}��� �O/s�U�w6na�hE*���l���G�>�A����(�aF;;���n�ʍb�Jؾ	w���)�-iʬ-1q'5���d�i=w<����b�U�����&`)"�(�����lB�>[���I��_i�q�+�OO�$B��^1xx8{�-R"�@ؐ[-�X��"�dh:Ӥ��e�l��LnU�]���\\�P��q!��k;& |�s��(%�r'@�ˍ��`�,�佰���Ԥ�pӃ�3҉Cd�#���D�㼎=��;�5%����i��֎~��e�X�?�% ��[�8���Y�[
�f�W��?����.6����oIV�֔WZ>xr׬_�_^,���Q�3`�lq/\�@�O��pe>� ��<F$�^�M�$-��j��*���j���]������-��'`���,w����C�G�p�._��Q���0Sdѐ�K�?�hu��+F�`:�Y�%��׌͵�0��:D8�����Yb_B�{��a� Ԯ��,m���*`�B�키xEI;�^�{py��H���Ό:�����|@D;�Z��������p��'xR	#.@�V&RP�0�Z�Rz�({?�f*�����ʟx	fo	c�� KF��	�(�7s_����
]f�ؿ��ov��n��Ŧ*k�l��\��H��>����!�Ųl�|��)��!�)Ѡ�s���9	�髼HZ��+՚mkHx�.�����Hq�Ժ�	�.�{,Bx[C���հi���d���p4St*E�J�Զ�U�E��Ŕ��F,��I��y.|�	KĸF�`/p���%��9+�eoȓ�8N���u�Jp�y	}�]�t*���xqA4�!����UJ#����
Fo�����Di>۫N�a�k��:L�A�{�VĨ,��4�?�`ߚ|�1�FwG��D�Y���ݲ�z�y�e~�W�b�3[�/��Cq�sz[0	(�?�`���q+�BƋ�Mb˳��e7�n�6�I�G���p�
<��qCK�wE�y�5�=IjjF�-!a��4�K�	�s	���p[Wo`���ɪ�cn��ҕ5L$�!��y=�5��0O}Vv0峰�[�"�����.q�3}�c���rm���եJ|�3T���Y6�'%�;U��p����]G���b�Rr��wB=����~y��)x!���fg*�`�8Q�7�* �-�']�Yn����f��'�����6��^�V�<�G.�Ӧu����U�T{N�SJ�o��[�
@��6�Q��!�u`0HXi�\����P:Qb�GЊ���=��?_�
>٫��a1�����T��UX��ߕO��}��97Z���źj@�����4����B܄a����xVb���D1���jl�6��0~�i�n��y�}���Z�p*��/y��VT%�����X$}��x�.�R�]��3�W	I�������5���rzM��ܲ���)�sC�ëR�#h̌4F�-���qͰ��F�e�V�]=�@%��O�7��A��c�Ⲓ��ԃv��P�S�9�	��+Y�l$�B���8g�g�:��4a�z�)�=���
�fw�����,9q-��Jy�!�Y��Q'�!ǩ�l�+��R�x������ �˭��JT>���m��`^M�H*��������k	C_�d�}���ۏ�P7�_���27����V���<~�WW��WT��6��`�wM{0e6b�/���gbm��\�~=ւ�AP���ђ����K�^˴T�P�K�2��#�+x֞�T��͇�m>�'�����R����
#���٨}O�aW2#B���&Q:�b���E~H��߹i��X[�"���̈P	mee�2%Z��(����@�]%�`�љk�G�bp�*<=�W[��U�V��1��ђp[����&�'��v��m�v��ړ(��	$��*͍t�|Y��S������>�A�hu�Q�+�3��D�����W"�21��s�O1��~]x�F�	�tn-!�:���� k뛈N�[O�C� ��R;u�Kt~m�n�
tb!.&�Tk�`+�u��/�1D[��S��Pdv�Я5�J#�G�>ل� /�Y�S�*���9+��|0Y 7��;��Q��]�i$��P1+�+���z�����s䲵�!�/j�"��Ğn���Yq�Fy���K�d*�,/ï	�9��6� >���p��V1F�����@��������qn_�<���q�:%��{���ǀn6(H�פ�͹u����C���U����J	b�%W����վ���{-Y��S�B�$�T.���?�6�Y�õ/�O��>�T���ß�X*��8�VȡBD�~�C߾^t��C�w#�G��[c0�)��wq��B�x��Yݞ���Ͼ�V�A��p겲��0�n�Ya�w�_�zM�6�Ք��B�m�� �4Ri�f#A�R� E��$�.����$�&�Xe�k�V��u���c���6�B�X�{�hmiY��f��?-����(�۾��Z
l��?o?~lqS�ge=�r�w7�L��ח�!륃L$D�ύ�}�'���o�?�k���� Lۗ��{�̮ÓmMʋ3yV�O��l��4�B��q��{�[ݒ�R��3�E8#n���m��P��pf�L?�@W	�;��Z%��eg�aj1�+;���}�^��
�	�������RAJD��.�����	䱔*-���I3ٿ��h0KD���oo˴��s�i���|�U�[�6��k����?P9�!�׺�i�'J�:7#���CI ۈ�8�3�V�hi����f<�z�:�g)�]�eW��?�Z�)�� �����'3������|�����"��s���g�'J�)�]{�=�v�Åeս��6�A(x����4��B(0�<T�aw�B�Z��{[����]z��8��L
 ��h���H�X�Fgp7�:a��+���v��0w��	�O!��BY�,������*�����, C�b��\�{�Z�|F�>4(�r`���.5|R��R��,D@�"�J�àX���6��`�b�t$	�	WO�>�x���drp!0_�^ J&PRU��'4�&7bȥ�֛.>GUL��DؼтB)5���&�P�	�X���n��ho���w]�Tw���Hz��
��`@}x���x�� 1y4����~�Ց���O�OѰ�h'���rA�X�Z���pڄ�O�B�6�����u3BI��������=2^�n���5�Y<�	!�c������o�8���.�{P��C���FU�y�VG)	-�x�j�Y��0�I(6��O?�#Sej��B'R/p願��lf�d�A�C���U��4�@���߸��O=����z�3[A߼�9Qp�*�;�A�3I���(e��_�Bn� R��z0<��^p�U	D<=P-B˶�`��\q�1{+���Vi�߃̿X[\ &�Y �$�z�6�rR�qDk�"��)Kn
�j�o�)ِa���`~����)/�W��$'�g��R<}n���{$s�X3Q�E@���g�R�s���,�"[6p =�2Q����Z�7���z���+dK�]n	?��hL/}��ȗ�X��pd%�=�Zr3Z�q���T�1�~�k�᭨2W�l/���^m֫#�����Ǯ�@U>x��	g�IL�u�(�L���>7Q(��f��J�^���:<Pu� �}ܚt�Ĕ^]�7�9�!ɯ����t�����#&�߰���烝���=����=nӛJ��O/p�(˩��Y��v��k�m{9pխ��ę�@���\��Ý�T����m�6���K'��c�	���E��
D��agja�BY��U��F�V���-���,~�`�)�aݏ��*�q� a�<4�[��U?ܜu�"O�L��$d���zq�&�&|
_q�s����	���_��tU��oh�Ֆ���_,3kuF.����D���g�y�GjPnQ�q�������/?��aFqf<����UN^��pųb��vK��ZZ�2�S���"��	n���gk h���Aſ�ר�ÏTcN�@jg9����O�P���0{��+6�pgs�"%)T�	�N����zr��oG܄��g�=?/��'���9���7&��.b\�#Ϊ�c �#��熇�N���o���"�ؒo��w�����S�m��m���lQ��[�E�H^��=3u�\:A��	ݔ�M�M7�����0)͝�rn��,
��{H �	-�8�_ ���Y7z~@Ϯ��q��a1��B/�l&��\���3���K�A��St���B@
yCR{��C
Š��jk����NPP#����d��R�h�,:pRx��s}Ŭ���O5Km���:���aw���3;�NG�}�	�tOP���/8OM�'�WY>���~Ni�4���;��9tf*�b��M�^���!8�%��_e*qzh
�����G~���������_����� /d�K
(������
�'���SR0�al5P�B�e���?A�doR㊭����*���5{S'i{���v0�/B�a�M�lǚ{MKn��4�8���`���O�k\�^#%x���x�j����ʾ!���[<y7o�.X�+���0�ژ�_�\ �#�S@&rÞ�9@޳��A�b.A�Vo��Z'������.�5�^0%�����EP���wO�,V��+'�Z���:6��v�e�l)w[z8�D�c�0��
�hg����0� ��˔������qe�ov½60���w�a��XE�ѷ��'O���V�|��_��Qf�ʙJC5���JUڨ�*�wQ�)%������D�y�.���,sm	�{n�bEF鿘���) 2�5"閆�}�z�!L��P?���;6p����ђ3(26�T�5:��ļ���H��ƅ%�H7S��T,^�y@j��~�j�D�A,o5L��\���0�d�Z$���j2hlb��X�O9T5��,�<k��%7�k�cbw�4G�>���  �U�:�����dw�9&�KF�ɩ�6iK�~Toq4�T{�c��Ai2���J�kR����Ĭ��t�~��H��R��J�3te��U8���$���^�M�Jk���;'SL{O���t	 ���+a� �^X�恇��y�!8�,f�hp���}D��>ܿ2(��%6zls�q):�TM$�QX�SRk1@b��,���qʶ�a�FXi��0��G�ݢ#p��^�X��2�J�t$�U� �ѧϭ!��u�G��8X
o �v�}��'	�.�v2y�#V/�n�,j���B=��5Ǣ��v*M�ͅ����ډY���� �u�%�������'���JXƒ��}�F$n�������$��ɵ,/��n�_+�� o:��1��3��k���XM�P���o#�(\����+�.?�:N@��,!\�2\,w2��@�4���/�����{�)�i�%�k�8H b/ѡ�i����M��L:|۩-��ܸ#;��$Zum2gt�Ǚ�{�k�6�G�t��T��p�*W�C�^x���3�[�n�m��l5��8a�c+h�#RJ���G׳�������
���"΀��թQ���`b������7��<YV�V-g;�~�.(�
��+�Vy��ꞌ�����S3<�k>�#���P������E���x>$�|J)/ A���>�e�^)6��茐��j�{C�����e5��"q+G�b>c�`�/g����ը��	,�?�~�G���⿚�X;��Z�������t��.�8=�SL�tON��Ƥ_b}y�"���܊��4pa��8�Q[�Y*�k�$B񧛂��ٱ�1�����g�����K��d���Qj�&b�U1݊f��z��P�K����cw�9��@��������z��˴�&Wm��X�ʣO�����-�P���/K%'��U��׃p����1�}��M��
K�y�oE��@��9]3K�Y�&�E��X��1����D�:_d��b�	
1d8!�}y>f��3D`F"�C �D�߱��F���RNV}�u�:es�'�|�����בD�Zb)oO[
7�������&r��ޱ�m;�J-È�aG�s��N�S�8F���հ�v�#,�2lM����?���sc\�7��֘K�<
e<y�|}X^�+�%̹.uy~�zZ6��Q��/V��>ع;i��:�� ���l�O5!e׀H��� L-`T����@�����];�Q�=�Ɍ�3�):+j��������/5j���("d%��iO�
k�4��zt2s��V��:�3:�U��#p��򨇛t�ܕ��w��/E��b�\v�n<�,�ٴ���o�#$
�jmV]4L�Z1���RX�ksA��4>E��.aI	8�M�/�E�w���=�"��5�JSQ���{�#a�K��v+	�(Vݒ��	��RfO-tm����E͑�4Q��3a�о�к�!�O�Z���=����tjٻ��K#�	k@�=����M�;�c�m�5���>�(�Ԟ�jI@�UKJ+}p�1��)J�E֕	t��4�:�eD��?�|��5�&�T`�̽�r���IT�*����N:��^*C_D�%ļM��A��"��gJ�Pia�r�n7ucIHҖ A�e=oŴj�˒C�L�_��\�T߷�Tg\Zч����Y��W��]y@�b��8bR��9�.����O��S�3 S�����z"�K�zI\�,�����
�X�Ǐ�>�L�A׏�,��AX��I�V��p���N����˖:�Mݬ��幨�T�o�g��Շ}(?TF]�K�!V����{i|B]�^���Vn]h�Y��y"q	V�q� ��KT���qr�I4��f�#�6'���Ս����c����p�i� Ȍ�B-��˽���2׋*�����5����20�H�5^��P�7�P�$0u�~	�[&7�b9�sk|��a?ӕ�����e��p��D��A�fր�xթH�P���]�
[����x����	�|	KYq!�&�iщ@Xؚ����#6��Al�pO����9�^oyT��l_��������?MIO^	R8�aLV��h���� }H*��b]Vܭ�yCPH7�'y�#�B�@,I#��f*�Ǫf7Q���|DI�T�FD#(l�k�署��f� W+&����!!��@E
9J���@^S�钕Ez�����+X�t��O�B�	�ػ:hQ�M֎X��(��z�g�rìyH�Pw�KE��1�T����jr�z`���'��*��T'T7%��K��ǅ� ���	�����>'3�,�G		%ǥ��5a��6`5i�_^7��j���7��v��g��{h����*;<�7��b�(�*��Vd��d7Nf��Z}�/>�N����~�x��m��_h!)�6��%���#Os�@㣹�؆�V���zz�qH�wL�����p]���V��J�5��-
l����Q�`�1tk�
�G�-O]�� Bq%����zo�6l5)�uxD��Y�/:t�
���:�j<~K��~v�Y6�OZ�ϼ��b �� ն�˾ur���W�[��i���U�?3���79ɨ�{�5C�}ko|u���p���V��S�Ë24f�f�������f������$���T�`����|��-K��� 1�&��|�E�>$��hh,�w{�D��W��
����gNW{�����8&%�H��A�&���&���牂R%(V��6�Z�`Q:�M� �W�b������2Ijߒmso�x!]�����D�V�!�o�5e���G-�6�Ҍ���@�6D�?�[	*xpw��|j��h��F���M^_AC�0�����إ��HCh=�7[��7|�E�18��V2�7c\��C���k�Ёd9c�o�,����������nz��Com�����<��W ���>j4�Рp�YuѪ8"D�H{MU|a��K�k��)��F�M�&]��o���[�o>j��x-* ���-#nx�����`�9!k�$�?WK����<��{ل��!�Com�ݥ���f]o=���v9UY@��&��s�L�!�k�R�I��#����R��]��m�X� x��oL�t����a����A��Щ�
NH�˫��"���M���6�
�Q��a���;��Q��}�1D&�?�"#R��v����	�����<��q���1�z,�3g���C&�+Ǣ$30�>�L/��h3"�Ta	"����#��I��j�?�O��Fs��_ՏX�|� �?X��,>�g��d�U���1,7tИ��}��\�,uB�]�w*�`�f`�7T�ش3NL{�A�wdD��f�=5��Q��Ք����'��=^����R�k��!t���.��N�uǲ���9(mm�Y[쳅���y'[,�����-9DGL	iH���S���4�
�>��S=VJ��amArz���`��.!6`ڼd�zW�3���UT4T�a'[�j���.RMGZ�;����݉��hW��*�W�`E�ܓH�#q�`B�DC&���C����a�����Z��FESŤ�!����ݞ�"nw1ъ��@U�r�����v�� ĺ��q��jt'�lK)(�a��p�K6���PC`��4V\� �����E��Q�?^������%8��(�n�Hl��N���vi�+��4h�>�8�'���I���׺("��яu+0W2�a�i�����>U��9V���`�F���Řѝ=�����w��A��u�#&�S�(ؿu|k?%����=B[e�5lJ V`�!�'��Q�t2<�h@����V���.�~��u"씳᎑�um9����=F��VР ?�����I-j��zb�1ߌ�W؄+Z��g��%[Uw霊�+�+�fR>��l������>�>���A������\&�n�.W}��ci�a��zK*�׶� �2`��X�.LX ��i���R�c�C��Mya����0	�n�k6*�3v��Z��9<�etkv�S����/S��l�ɶ�t:u��#֗l�>��� 9��}�pρ^����	�E(�2	H����Cx���;��1���7{[}��2!�$�s�VY0V ���kEO �r���q!�yj���" 8|䳘g��O<gN�������P?Td4���,F��x��͉��a@V�o_V�xľ`�����E䪵k�`d��kk,�/��o��͐ ��H�en�5����4�U��z����aD,�%�Ve����<��m��|�$L3����sK��i�"$��Ү�d���H�߯O��Ѻ��ƻ��8 �Hk:�nRF� 8a_�����B�#JL;�'p�fi�����&��*C�[dr.F�)�z�L������VGL�O�o,#��~6,��:-5dQ�\p�k�@��+�150d^�@���kWɂ�=��ҩw5T�,��֌�\} g���k+��
�cr$�x?b�}GͼQC�4�ˈ�|�ۆ�2u2�h����f��D>4��>qag/���n����P��YL����bĢ3:�+��j�2Tx���6\�d<�Ixpzێ�D�x�EtNhc�1��t�P		�q��k�S�[�'�}\��[�{�x��n���NX�m��3JK#��7�[��M�]g��NST�ۗ�M%�e�J�����rL���Tt�h�Y����x0g���
�yI_��c�'U��?�!K��y�������j
�IRl_J�j�h.A?��� �!�7k�j�}���Q �}H���^{@,��)�R��hc�,U~��"�� дg�C,`���0������@�K]ֶV��̂ ���4��%ա-S��\�S���!=�e����c�8��Ͱ ���*��?��5 �R���s��D�
�t�<6��Z�":��=p���0^"��~�V��e[���&T��̺&��g�.
e��"��{�	�m(sL�|�4�sQ�}aH��� T�4��j�1-	&��'�*���d,�n���R��H�٦�]�!���L2҆���Z���8n�Q(�v�}(�C��ԗ"(u-���*�Ao��5�5���&j��1
���; ۰�atZ��>A|�YGn�Blֆ
�*1�5�� �Bl��7�;c���v"�ht���9�v�x�{�����eU��*M�϶��*p�\ݝ�����U۪כ5��-PA�<�Aѱ��k��GN]�忣h��N�|����]Z�98��#`�F63<0ǭt�Z2���Dd��\QӉpȺ�N��GÒ��xf^�b����'v�g��m(�?����QtDx1��xl�3;�s�+�rE^�&�KTA�(�Z�$���0$u�?k��.�e����C�ɸ�d��R$ 8{�p� +n����������io�{WC�Y�K�%o�c�A�5�� 	�*�#�t���)�q�Th�<P� qb](M�e��w�S9	����[���񑀌Ыi6P���A�A���U��r�w���y챙2k$����հ���(G�V�7���M��ɔ8N�"'3��e�-A�����L�,��"y��(1�7S��?}�G;�����;Tl�ZIX�k��5�<V����ϟ��ꀚMCj�~��r�9�4�\�bH����$+�Z���X�7�-�޵�:p?�D�)�=v���e/�'^a��Ǽ#���l�1|�� %�\�8�$��V��H4|�L�;Q�<=���O}^[��)엜9[,禕z2q�
����e�PWQW<��K�������ݝm��;J��<�!�­��9*
�y����kO4�����ؕ����2'�`��DH�-��!jm(Q�N�Ba,�̖�8��+x`���n��m�Ϙi��^\��ތ����}�Q=U�<ӷ+'�J���('-9r4��X�x8����"e#P̉9Z�I[�w ,{�;�9��P��?]���{�Mv�<�v9u���J�Mt���k3��Ơ��;qa���,S}��+�Y��"@r"=�ʢÓ�OG{�Z߀ac����G���y�W�O�U����Զm�g���������9� �6�� )z�Y�q+l��IW�V��r��<$(J�~FC��)�h�\$d�C�"0�X�P� e����^�1v1��oD��KT��4��e�7�~͵!?��?��R�_�n�7����a]�
ɀ���%�a^$a%�_N�N5&VW:�3��+�G6SM��,g<k>��bC˭�
�>g�£�X@��<�o-�F��^����N��5k�U�Dz��L[ @ѽ9(3LY��{�� $���f��O���Nw[Z�4����cy>_��W�9aͷxp���q�kd+��O��	��4�vb��=�uڋ����%"���= rI�0:�;4�/j:$/L#c��NB6�o-I��E�f���{���0�T����b��b��J�Ůǘ��n���Lt���Z��8U�FF+��Go@��x=�֗k(��$�t��SMl��PM��9��N�Y�i�<��Lt:��.�:a1m�����y�­�F]���e�7�	K���ʅp�����'>K�"V+��C���%��8pEI,t#���dg��L7˧9m������=�d����I=u�=2�Ma�Np�r�;�eUn��$ ��w�l�e�s�>O"DI�&��T��m����ʅT
h�#;�;��}v��A���5�l�B	8T,iԾ�ɬ�*"�B�� �G]	-�d_��r���_w��Ʈ|5�}$`Uf�+9Z)7���C��K坏y�l��R�%�H]I���Q)dv?sL������F�h��s+g�Jp�"+Y�T��/����Sp��G�1a;��U"w{�ǖ|���?���Jꇢ�P�����4 X5�����&7#�e�_v�g��RBþ�ŀ�Y9#2�픶���U�ӏ�c���ӕө�uH=�/!"��P�����@��#H�fSD�S�K��+����p����K���F�LG�͹��V_�(�Sl�$U�I9 U��x���}7��[�2��٦�>`wP��/�P�u"Th�^ە�4#%4�U��ݒ���J�h1��$7l�lI)�����˖?GʕV������:��(��S�<���EҮ��g�,�t���[����6݊�q[xJ����Xy��ʕ�3�k��L�Ӣ���+π�	�)Q�^�@6���9u�=��.�E���M��#S����6��l�ui�CH,pq�b}L�s���
����.)�~���qj�l>���$�yz�^rl�: ���}n���Z���y3z�ң�;)]�|�r��4{�st��[�g�]��6tez}/�o3�u�#
�M�܉՛�C���8�b3��I�$#��Վ���ݖ��i��@m�(s�n����a,O¯����G�p2۵��|���cF��gc����~��S�Ɩj 0�s���X�h�^���+%������B�M^���9ᙒ>�ۗ3