��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a�����{������#��j��{��	?+�g��-��"XSʌb������;�b���/��.v���9�Cl(�l-i���C�٣ϑ��c�P(?U	w^���"����Y��j�L9-(r�i�{�߶Y>�&�E?��;/�\Te ;s�f�0�����[���t`Z�FE���8)(�v�?!�A�ߪ�"Z���Ǌ�_�����H�V�jVT�f��?[U膩P���8�K{`����X�$�	ʑ5\�0j��}S�߁:�^nP�+IL]�lnUSV=h\<;w�������$%K��]��9����f}�����t�|�2��iu�1�V���,�� �F�,���Ԯ������Vl�R8�r;3�U��Sz���C�X��%�l��n�]�]������V���:��\�߸��TS�f�XG
B� �Al����W�6���}��])��d�#7p�@���c5śdߩ�X�B��`x��N����{�>f���K��I`�Nc��|��<�� ��d�
�!�p�D��w�]7-޷6��[��e�Ya�xN��ẗ�� �G|��Y-�>�����?TFB�Qy�g���Q�5�5� h&>w�����8¦}0;�8�$��.���4r7��\����e!���E���$�t�>Ȗ��g�[�U]���ѭ���*��������Y�ā��o6(I�.�0Lߚ��<�vh�2��>��z�D/�������E�(`������1Ju>`�s�Ks��ˇ��6z:�JP]m�W���78O�B��-EϢC�@=�1hV��rZ��(/��R�S��+�<l''�$m����K��F�@e��F��FSO��f�4F�~�^e��!A���r���(�sS�7�!�j�x��2i��5&���Ym9�G5>"hP��|�;���!�m���ȩZ���_�_�l+�u������1\��~R�3v웁��B�w��f�:l�1SEI��}��Z�����o���EIS�@F���g��\�V���ՁD���\�t�^���I��+J��{Sy�4d��u�5�?�7�,����y��}}�&R���Z	~}F�O�Ԋ��k��C�T�c�g	��z��O��.��"/yZ�ƍ�1�k5�t9�h��殊7�#q����O>�WhHP��p���~���̲�����y(Q)�[��ߵ��$��d���Iu�{(���X4�w���n*���]�,���;p�'��2�� r��赢</�t�ZTT����dP
9POn$!�