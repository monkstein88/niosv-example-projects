// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
hc68kPBMtxLuG8NsRFBu/UHC0f4gkZBw54DW6Mh1vyggzNC8MV6mbWLW4JmMYDp3LPFYUCGdYREc
Xx3AC/Kmw4/JKVbd4v4shUTG5mdRPuVPzJwubUHk0naK+JALI/n51XeJ/3HrCXZ3q5EBp+psSjG+
8yp9xo6+bq0ANHynfYMl8et/PveR4JPXFXE8M0C65oJ5s1KQqooqeN+D+BgsZPkmxeoHJUDuHywg
GgPPKazZ+Aaszx+RM068R4BX0PZx1YEQiX9vzlAQXeVY4rB1lkiPfYEgmI6EWd62mtEWNhH5Bhox
zTqltWSpKbNX4ZZpqBEHlD+4hLmXzLw1LjVciA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22176)
91luD8yUQuHcwUSkrxzc/V+GUBYJrMiE0NML4D1aNNGnD6/shoMSRZdUHPwbTm24EUlTP5aDxGVY
RX8HoNRe2TrAGeeZFYtNR5NtxCpeY7FA54eEAy/jkYWpz1V0x/bPr8F793gR0zVFnroHcApJ6MWq
LSNqKGrd7mi9TRPLIyqkGei0z2jKqQ8HZ/6Qc4V0sO81NJAtKnbYNWK0Ic/O/n2NLAbCswDkAqVp
7tg4Ldz3+sygZC6ID075W/wnqGOWdeRq4sx/f/O96SDcfHfQYvB2O02vQWvNNI6glV4Bgv0gIgJc
7pMSiH5EAW4+5s53HN8Tbr4TW8zp8JRxBuXtc74H5aOlLfBlgKIir3mdwBXok+aZ+/otousUw9df
UeaqYJ6HeqVHYMlFckZs1epbmJQDrK0lNn7JCXBl/GpwQMGgi711dlo1/vs199zepuai4ipJltIY
KBoS7Bihsbl+cVPniDHyxS9DJgE88WYwk5q2Q2kDG5uGk2yAkE6BjMb9sgQr2p/7UHkz9qjXkw3B
qsA7CxicFHsVDdmpVJSk6gZgcDrEwgOdgmkRw8OgkMzQh+WYJQMWhdGEDLK0FweW1qtJWcWCV/B3
fkfNqNi4gy422cOD4/uEnyRvyaaM40V3JjyrbDgwLMdtlUFHwrY0NEqHxkXjWCZ+H0ifwOjQ4NsG
H/LFEvR/KhrQGrLOlAqHZFWU6qRjcquVbkdxLC9HjlunCq/5sl7xvY8OOshmlaXv1qPqAkbKpQzQ
XyGW2aJDAVKCu2QiQ6beucH6fwml1Skr5HaklXm2BfgHF+OGFJJuR7J+WCkwPgdgeLfaqcq+mMWX
WO69n1SHqneePFIA4V+vohvSo7T31Gltpe3ge1f+7zEto73gORFL4Umh08HuhtVC0mbEesmLgiZW
6iSYY5rwle2bCpIGY46Et7snhSJhu9a2eyGgdBKW8/8xQRDhVENyV/nxuySDt3cJS4nn3GunWULa
hvjboGsAuCBbSxmeeaJ2R6Q9Lg2Ovj3kHy6zuboPxpIg2vY4XwlFV3hkMnPkoHMjuTBdgdA3oApW
zN73mdeGHd8j+JqTpiqG7rUrPz2cmFglRUv/6YjMaL5AdT+FJsywYxBbk+EHuhbkItoRn56ai1QN
nV6t7GJz3Z6WyhfCa+IFvCexQ/zcfTDAYnW5bDq03ext0KYCOmnXt76Fr9Nin68i/WRe6NwzoSUg
Ay5FYMFhnL3hOpY+5cb7MA/YQxktCHszl1Sn9kqHAnjLuSytkG6KNHbQE8pj87Y/8yvo2sweyFHV
40j7nmlzA8aYozzZivUx072yvRuDhs7Z385EWI9PidV4rz357/etZQ1XuoRZeUR9ZNwoJcGfiCj4
4NkrATUykag1doGp4fP4+VKvUBH7pb4JWAL9gIdidskYs5YTiYWepHdnf5+Tte6sdy5YDmLTInxc
YfzEP1tm33USPlF2Oj62Vk671mZMKGTeWOzPb0oTS04TYn3KB+ORW20maiMN9EfUhyFA5AJqFcoz
jF6bZOnrxdcbpe+W5Foey8/XKb5ejIGLDGh2CDE0nAVoAdEzdLGmmJ/itjxJI1hYVOFaxqGDV16F
tm1RJrF0aJJJSkQc2llYRdx7GAgm40fJ+sPsxqmkRkmH5dnll2DmQCtTSzEGJFkcz/HAtOC7+K1C
TyMw1XqPfR9D59Ovy0IzltI/u2kyIgHBXaLlRSmOTMGanwT4LbOpmiBgPpx6USh0CqPjHiESdmV9
imiameOWJfUw9c5HKvVFIT73AbLKSFx/R8jLBthCeUN9sE53dvMBYGsJ0x0WKLmKdeELUk3HNW7J
sjwr6szih7+bnrtrftaL49G77bvQzZic2CvuQ2FjYyRq4tSQLN507DRpBwUbZUDhyrWLjMgXtgC/
UvOii9vBf3b0TyKhRdi5DZle7w+SAaK6W5rc8Sm787pjV7nEWTNZX5yBjuDtdFqGOO5cPA9qkhJC
z4o9gmWCah+JbNIdNIVl/Sl35q4R8kyrkzp0Y3M81f9ltjQIul41J5LNlrnLHnZ7Mtf+Yzsm84Mz
uN1eGKXB3MG8ewlUEhT/db+JlMp/f49/vOpxQDubOMaPgQBNKb9UqQA6dM2kbLCVtSziyTxsUrNu
PgZ4tCaPFV/gNlNc9vJdJjABTqm9rpsonMyl9uAJH90eJA+mvzgTCK/ZZbtA874ehpRQaJ0kZTc2
VnGW2PR6X0CT/iImdTqTX6EXtm9rYl7HshYKLn06/ZRjfIkV96j5k/go0d8mZ8yjAw6uDzX8pvq/
CwHgvkOET7Pepb0v/Q5ChLtoBxOl43HmBkgCBIU1xdaGD+/EdAqk8/GJE0TsiuUG9nTLfr+uJ1EN
+3dNy4zhBLQwzFWAnFXCJxFD9FMDwQ+EixA56TAd/pW+i/3OJgu56JgmDYjAp8i7Y66RkFrqD6OH
ytddaeo24upbPCVtFCTO3bM7I3Wt8eI+XY/1stePM3ZVry8LN/5cP9MRCNjh+m8Cpn5C9pBSPGBS
0bERW/777mxdVeiZH8RHhhwkjtCUOTJtdkUVKZwF883JnUryvcERC0vaxHph1qzHksV3h7CUQa6/
MOg7Nnf0GWAnCY8+9fgAwfnuDjAjayHzuFMCvmSh+dPlXtlV6WDDJBXgrpWAVw8SxIseaL9aJvCC
ZMFg/Fq1aIwW4uX4DK5TQIn3ZNJGMyLuqM9Jf+Ll3W2HjLHwVQgC30XVfgI+v8yRv0nOrOvT1iP3
3vzd5PfAESlKzwq2ddyyUjMWjmw+WFgCS+NNhiaNxoQbBkrWKdWjpFDBN4FXMHEHuVqK+eVDTf/s
ho+g3gvquGkMiGCkH1Ef0JuUwzF/B8MVw3ZxAfnJY7l/VM95shbf+DXEGN+dQB05JBQaKcDgVVsD
9jRWVTWgy+xKhEibGTju300qs8S71MwEbnsr2AKhx70MLr6qDca3mKIhe3QezyqYPkxzG/aEHZu8
RRX4YCVsKKnq6+tT8JEa7k2tSxgIeI6jHPSHNjLyZ0RBoAsgcgiowtntlf4fLfRtdXUHXgJi7SuA
VtEifqmc9F1K3vKt3UWAD2rEPjO3t/NxFvkibprjFb2pp0p8QhAji3g01i+iGCnsPLVxSFAZAPi1
+nuicEBmtv+PoxgVDDhJAkt908uNFc2tCLrHCsE0vZQNTV3cAnng0y2OulPZcPsAynNqKUnPORmI
UB3S8fmZaegrd0Iw+5QuBHg5UHDot+uFF/EFE5Memp2bP9eFU3A2MfXOpQg804tgNyLEWTT5mF2H
h16BNDT2SPUaJ/DyZOusfSM/D+y4LK2jjk9cAwiHHuzp9/3HccPlB0a/dLXqbzHjK7gV2TVG5uE/
cR3Ix5XFVQ06aJ39BWaXB8kvsbtdmHpZV54XuoJ1QKLfz0A9oon8XdwjcaAU6epDn8uHMT1flNmW
vRTOqucv8B1qlGCcJFINumC5N0+2cIZk6iLi6aCA9d8SjxNSQngJILPd71KT+KoWsTsF6aJtzymf
yWVqooR0c8/sYejvKn/deXnox2C0pXSBKqZW+kSH6qZcde0TQlKk+mlSq3LV37u3skqQ2daFuB2j
gfhY7QAyZJim3Oo8bT7obCA6T0VCvOMjSK1KXcvDoWQ36J4MeuwB8zBpGY5+7YV9WOUGW20nO75T
6OjeqPu99cMCfItJ2ykC/uJNyqhxrqdnX3EFSYEWT1HJXFNskG9VPdcmiSnlAT+ijV5u9+D79Wf+
eKOIEYzxyeIF9YOlcmcEVt/4iw//oQCKTttUZWT3Vuyaud0Q2l//PS0LaPnC+2CsCbDwEewe9fhZ
3JWKt68kijdTXkys4NZdNGR+LG6RN/64FZ4Or3Vodgwr35BNOG/LQDSRCOsCBsD7ec7IHhpx6ZwQ
STNDu6Yqh37QdzdCB9Pw0M2gxvr7Titl/S0IBRlk8O2HRR0jOScpXpQjdNGJt/NZUM1lBEedeeHQ
yukfzPH5wcBfQa6xVdtx0BnsXObbxvEgd1Bgkoj4Vy2jQZwVOeWf9iXiivnMYP7qukakb0uqSMFh
+oHuaZRb/phdiwPtrboXiam/+9wIytPsyTEYRsMjSujdHxNQeFQvQDgsYOh99V1+620CyBbk+pE+
wuNpvO06ILYrgVN9H9UKy5pWIEg82tA/kJihS/TAZPrBUC1cuo+bFQUpzfpCbD4dXlEiypw+DU9h
l/A++zZNG+XA2I2OVwq8fdIO3tsekFtSvlXW7LYt+CaiHSzKVGaIawYahVKQ3mudq+S+j8lXLto9
J16bim4ODgX9e4qsQBM7OmVsJHg7/gyzR5oIs6XjgxCoSRsTfu1iKx3RBfbOHfEUPHSl7Es4LCm4
doQcfLYgu3NKnvGATHMCC2NBfd3KLZcxSbOFYX+95lJmI/EeJ8eTleywkW7nKzdPOc3NOMtP2h1k
kOiAsC0etQpUsVDEie4WfGZ1pRnm6jv//liW6ALkMwYD3HlOGrvpHkxN7XyPyUnyXUCZW1gq71Fr
jd68jneuaM5LM0Otc4/PMVMnIJUXZLOIMlX2CL+oeAVkcQ8GsaaDiAjuGL4ZsGqPwNGR7aaopLqp
UsPx5+QQ0EiyiOMjR9wJXe0lCDunupRCEOrJlkJ7hW8DG8BrcQhu+3wDyFcGcz3Tl7KhMkfqvEaN
8D+Hm9Z+EbwauJ8xTSTMP3RLXqunwqbeFJjGw7FArPaunz2lzoGw0aLi0hNQD6T5gk9ybkWKjETQ
TX1IR9X+zfCuwQfDhp7OoZYN7TVP+XrPmd0vdP3MvbVs5HjWGsHsdTDTQrgNXxMZTkQvjd7evduT
7DZQ52OsGC0cUMgFxzLL5j26yM2+9A0CLMBv5tx98woo0OhpntSNFMTPdNh6C+uNYIcz9oMxFI5o
moFqc2Nx/Otzd9PwCXduJZq75HD+JTmL/yK/Bk9xbwDKSIQMm9eEgqX1SLmHfOLxnXnvILGvsISe
HNLwJFh67jIhf5WsFGhuF2v6ffRDASFLvSWi/9b8xuZjXfi+hLVOjNRVNQnckoQwI2TgxWH2m0X9
1HD4i96qiLH8wOnF9SqYHv7QOPROXLJakr7h2DJq2W5VJGWTBqeUudaKbwRMKqRaGv3vdiSpD+Qz
ypVGWxjJyO7V2bWraCGIXVzcixidZ1RrcCdqSSH1wUdqpk1GVyOt8AyMAz4oHBAOI/LwHrWLUyGl
LWG2nI6pwnDbRT9SxVHWX5Nobh0RZNsW9bZp/1kqVqRFFMMhfSL/aUBOGL4WlJZTFJs4WUxOphr8
jkTt2HZQNsWxXyr+I20pL5/jZM5AMSbTF8/W/6ijha9T8U7Hb8+KiS3jWH2dqkaXEw+u3dvRn+7n
58dTiC3dzUQXHqhByCE+DTX0eN+VxpLFEbj4w1OCIjlRXvp3a2oVW1GN1FdWb5Vdzs7Y1IxxTevL
F1M5Jzw8kpGBIPOpIiwPD3Df9AnRNRjv/U7qyAxOCZ4yla2LQSLBbiiojyETpzlEgQ1vne9xA8Ju
8oIK7x6KPwRCPFQOtP8lbkPVAfnMveQNIxNp4puu+kQDuIaFlp0P9sBN2F8wJgCeo9Wlp+99W6Zt
tqedDm5iRs9CRlfouBwMuDlsR+xEyMz+V/dG5AFlRUKah9gmCQDoUoh1I8CGd1C8v0YAIxF462S8
vnWhLEoUmv4f0ShJWE9EOCdL0ZrqCU5oKSLiqKwjaOD4h8eOKk2rtNK5kGh3lAeQ1A9Ozlz7dLtO
3dMRiMpVm2zG9Y0TaO8x7BSpN7Mu1NMsYKIPvxfhbDHF2W2sCXL71+1VUOrUyfiFc7DkKqZ4eTuY
dpdk0ATQs6p1w7O9iN6NECWJvj7Tx+YkyZ5nsFrSogvxKOZ7db+Ah7GYJDzndR0XaRoC+0FaVX/N
kWnapd/amoIYHPX03lZNIaZD1m/bswzWdX6TrUdbFh6VIt4WYf1/IXDZ2MoPQBsMEXYY9A6OQo+5
IqyxciXddlKQROIzq1dmhCvGdtan+a/6r9q4U+n7UrvE7dgzjao+/gAKpj6HFsYkdGLrRqV1kE85
JZovlsNxj8IidkHqSSeanL925aEVn3kF5KtxSY3dJ5zjIFervnmnQoIelh+jWCPrPax8oQIDQtKs
gY2y03jEP/PfPUtJMaoEALokD06mHQ8zkzlQAvwF1Bf0MdnvMSWsT3l+hwmLi6jfVCYqwiLTYrmU
cDGpV/QtWp26+wT6YEYFz2u+OXLK/s9ufKzQwGHPe09BYZvIus5TFe7YlrssRlBfASAr6Iq5hlVI
AwRWqdOt+yTYig969Xef3/XjdKTj1my2EnFNdX8Jn0gWQYqgffOPohMclbfr3Z+Aie9x2N4yP0j8
topcPt4A3toBQ8olRvUf3ZJML2sxBMXD/Luj6GIfTZ8zPZKvieKtmD8KU6mSXkrBjIuwp1y2cuy7
XzaypYOL8L08bnzgeRaz5Dy2GKD2Q8TD99xf7AK4cBVlqueV1aGHWOW6vZ3ycg/c0kmT+bfos41P
oUAwN2hZnkuE7xs26llL1A+yECh4DgOf9wqipFs/N+sOe8QDLoK1AYFlE5mGle5ihdYpbRKNHQZ1
Xw+VdCUsvKOl7+03+C7mSS9uOtegSkGbwrxF0WDXXhVCWX3RmYOpxKX2qWZ8ozs+mqYrn0vKMPZ/
/z4hH+tVTdGLrdwSdvcuFSrQZYmRFEJeOlB3H5Y8Hbv86zvivjvDMnca4tRM+zzYbvdxqIud0BLO
PX9gf6T9mnQdmgerr1HtdoFDSNPNGH4NvtoG+AHjyUIl5r8CPJ6XCVA1rIUJHKVgpyMJR/1wBy2G
AkjHi6/j03+aCQHpwhPhNDya6TWQrO4Oqbio3UzoEkn1vFyivSSpNOqCCPv+IlCjS/8Gu9xMm0yC
6gLZq97HE6tJTFdZ/ziZFCLnjevNTA6lG9K2/IDcG+fDPKxB/QVo+ZNG+n4u8gDtELLgQifiscXp
6B2kERNo182EwiXGa2Inxk6zo8giSH6KtoBinJ8iWqmivqBXGesQ7gGZYEEtWIobLTVkTZhRxdkY
ZIyuMAqJTfL9IQdtdHCXEEitrmBHZkQ9kd08udzpE2snZEUcPErPfSAKHwBjrjJ/c22JjORZr/Rm
J+wUusvnLuoa/ZH+Pp4oRh/j2y9RQqaELRKzfPiNWLFnZRL8qtIeCgCKMC/8RyUlBdvJfU0K4tlr
nPko9FFu7nWMnkS6xymFSexLIPCKPnns9MoiiEHd8uyioyqo8Y2TpqaIS5s/Ua4l3cFZ/RhwJEy3
TNvRno5456jSj7UBpMTqPKzZYKiB5QwR5ETJzJA7sa07fgqA75P1JLIz8mUb8V4O6o1wzT741Qr4
hZVjRrhQMwnLmvV/u33v2tPTdQhtF7Gxki1E0RJ/ijURP2vbK5HgiBbeoDx1qjdx9BRTKdpMVyki
mhSdoinOuA017cbK86TCz5bUt7zhDAE5KwdVMMF1GsJrM/FKubNZwtPIW0AYlQbBPdwSaDMroG4/
eNxWzPdhQzp3SKT3gckZaSpC2676PFTwjDO67OUqYintJ0UoGb+I7hCdIjQ3mz9VQRG6DiJHpZ8K
p65Ltw/LPth15ckTqwW0jenLmSK86SMyNVsRBipaiMWC7mqEURAzuCF6vaC0yO7manyV1iYb022e
NUPKHkSjnJXxTDydpS9Ac/iD6IFcTg3lFhgP4ZVaBHwTkcj+2sL7j1NYVH5BoNPb0HyHBaK8o5t3
DcPz3tsJOR/EUu6jm8qk6892rk+7d4AutHa66PpHLfByQukFQ86zITnpNTTNL1X154CRIvZ6zbGw
Wn4/mPFQRFtgHn+qkvMzKvNjgCzkh1VvpEajZM1FGR7raQ9JSgsdPQinxnq1jwXwmZZLTgblZaYx
67AQLZbJ1ODFDIomo0BG5pfNp2tqozyYy4KoyHm/7bf7MTy9C9qCbfk0u8bFxi3MMckacCgpWK+L
yn4zirh9kjg0GAHxUHCNHb7cdh+hU7wcV2SWtUwtAG8FSh3LZURnRUqX5MLLES8FFEA8ESIBBCFu
5DCmy9WLyJCwFwcYIDOE5RXNhFxejuhL2pz31H7Dy64GYrAYiMQ7BXSUDg1kSRH/hxWM8iV+n1Nz
2gjSsfvHw+dCjyHOxCzb4Vvkl9F/fe9iqCsy0F4JaiIsOp5dbioBgR8SDdiOBWj2SN8GJV4ai5mR
V3kifjGCpUo+POSoGVDNrYKWlpNg8mmrv96d1350PqjS2hLl3sjXnJjaxOEZ7VSanY82nIY4Mq0O
Swp7oIm2bDxXfyjaPhqOmnp0k1suMYfBDp2kvdp0VqMJgT5qn5CsTURt1M4mgBh84n6cNoZ5GsQt
XqtNkLifjSX+7isWMbuoGL5HULhjLj+QLoeX4JzaVUFW3yGWTKkTzE+z8uG2XkF0EDZLjpsXS79S
AzAlV05LRAdUdGT8Fpb6M8t/cuwHnpHp2WQn9cx96ydy3+ZfSeJmkT2TjkJc9T0x/iT1Df7UBpMo
DH+QlGlezWbuHZkt2e7Vs6YWiJevoatPyObhvYTlRbqVXnijjcsx1KY+/B+n62QSYInMrrx76XHa
ndknoh+HoPLyul1I8VmGaDvWP3AAtFAsE1gnIWL2+g6KzL05KKUvxXEqsXRQSn8l5RauC6mINNOP
g2pBQIdNyjjsauM3x7t0jH50jQp6MTfvnpMW1HzaWP7VFqbK7X6JxRIdSTFmi0y61gAJqn6lRB1+
GdfueN8uqfSVChFUCRlhve/HGslkrPMboI/xg0mG2Zw+kByApG39bbwCebvOVFxNDxsvmLY93+cg
h4Lxl4eitwww8xP2xPpZldmYxPHSHDqglpchdZTRn66KsidpiXZcgJb4qOFr6Jep3PjXObRtya+V
Co+D4aCJ4b7BwuiBmTKu9/3iwavMcRnfRGaz7RCyU3OPY+KPbRUfpdbMVP+ad9Be/3EJGIBNOgl0
dBLeeZRwMnifIBjkVbV4ZfTeZg+qJRvDoxzyGFCwd1H+dBTjVKiCaehX6srn4UN9V98hX2DqgNRN
xyFu2q83jhUAM5OGOlmbaE1XbHsyKJALE1YKRaJrN7vbMvTkugswOxIw1drM970uyMx96n44JRyI
LL2IjOm0KQo6zL7oIqMPuGASzmxAMYuhJVKxrtoh6uDBLgmo4Txv5vk4DPeyBmX3wqv4sOCSY2C9
pS5TERQ9TlUowoPIHAAW1ojnqK8oeOL8rbq9LBhUWFUN2COGzGbO4ssux6I1WGRcU/Uq8Sog6vVG
bOIbevO+T4jxVZoFWdvRSHrFbwcCQximfouTCwR5JYjfSMZhyoltTuXDkSTCUUof+dP9gNCa9l30
qdEX/NKEuBV8ByXDX4IxGjndik2cHQTWi82UCOFZhaZ3PeDYINfhQGDnUS9I41RzaYG5IuNJfZy3
/vLMwY2lLFLfzUieVow3qYt8jRQbmbTRpwaEaZMaq4OAvaM8zUkqGMXC5Jx5Z9CmKt/sufZnDeMt
HLVfuR5lK9mFPMScP/MHioQRrbX7TGiTHa3z6LNwpXDfzeY5CewOKfP4llxhaO7hqIao8/e6IITp
f8GPrsupbZk6HVuBKNHDyNjC+Q9dIgnvwv5pc3Aou8Bp+6dqtvvntmQACJs1QO9uVLRHORjqWp4R
U5nkL125U4jR6a8sjAHQXgvlb2YLQVtJ4HDwj9HEQDVOxH6L9ysJs4e+v3t3+764ODbm20i8kK0A
E3CDM98NTZ3d2wr5RlVvPJMu22DEk0JKrM1QOJPcugbBB1GeF+lvObUSHb239e8c/+yh3AnHjpaR
aGTus2/uMgYnEYC9JjjkVl1xWDmnyFKtWLrIFx5NZUXJdL9fB5x8X0tRqEyQh2TlrwUMxMNH7F6l
vGzgcVPJggYzcEI2aWLNK2Je3yEC7u+B8YbVYaAl+Vb8ZfPSKX7m4rq36X/NBPUJkti3AzhqxI+a
VIRR9GKjxCxT4wUzYC2GCgfORZsSFy05w9Ljm1yGe1dG0swkZiiuu9aBQelxC3KT/0t6rNm01nZn
2kEzBsohJ1bwKN6bbkXSzcos1PifjTpadepdxDHhhdy01XOic3EKPfZ/gBk+Mi9iqXSvEHmeK3A+
PE9Js5yVpDVE+r8qUB3ymHevARaIfhskhWDdUP7M9ykoHBqt1Nbx+4iwT8cKtLj03x96R9povgfn
R2jM3gDpkQSD6vdjfKX8R7rBQzDvfVA1zQxeDHuHpX/S3FZgSlAFIs+Qja1GdXPLwNvS1SpcioSJ
8FkkYaunJF9ZQsmXni6Ec8oZi3di14vKOg/Tcuy/V9s4bVHBSSOWiRg7mHf/1ULtWZdr9pAwUZaz
4HZZ8U2h4vOS1SbeQDre6nzH+Mo2PDwqN7B2qtocNDvwKWD0aobqww8Nokbyp4SGbUVuENVxghdb
wLZ4tpAhE4gYXcCrLWQBBwRzTdXaHKH6BKPScGDO2FhaLI8m57WkQEYQtTBLMDpBg3Nn08Nu/Bm7
QuWO24ndUTBHHr3RODhd8tT9eT/zOMf/gfEuJcZaJR+fwDxwNRHe+aDqwCKS7D76Rz4mUOGCiPRm
99AssUc5ghmIgFVaUGbkfpwznex+c7kIrhu9VnZaEJLhlo9MOLxifyUdp4uL1G9wJtX6kFxDXDmb
l/ldRD9j+aTbEvLMiueg44DC1zXUxuy3zv6xl+/kYCkNSucH6oeC0UA4H6oXh9pAiu5/Ll4lWR3G
11a9mrjvm79NFYOmSvjZU//TlexjdiyG8pmvynHoP8Afe9XmG0VNgjCyE1qgRoZGBhbclhBodW0O
49koh2FefKZMkZzRGzqSlkhs1RJIhh7PhPrIwfKm24GfSXLnB2cBjA2rHi4S4r1L/knBciehLUB3
cLVokKo7Lorjw6bbEoq5tWokVfquS0rE7/SlmD8pxyCc1c1gKLHHLwpn4yyEIYdFhMt+eF+18iuZ
gszsm3GSCgmw9Ir0BodnwmjEQMhzn09L/ltad++s75FbrWAmcadm/uSJgoKge0HYty/vaWrJ6uEk
uRKRcyg22dQw24Ingd56fAqqCuEBXE7YB0ExjpOtu6DLx8rIIt/yP13Yhi470P1VeRigyOPKFPaC
rLbKSNYdm06cEnWet1RRm1IRzP4kAbIou2V35imhyTaDndG2jG2QB32yIrBGlJIvRxKBOm0DKW7l
gqB8EJLol5Q1H/7h5VSBi/D+b/bXyhS2hslPmZztZb0pmJ+VFYlYiBpReuHXeMhZqRNIPDZnP6z6
pMC/Q2sGlds3nrJlcyJtiYgL9HdsSz1NKqCV5SHXo81b6Ag+f1qgVtbLAPRpHFgtfEMN4foAtCjD
Qdxc4RnvYcZOg3VRsuTZG3htaKxhb7T5PL5OTi5u29bI062cgamPGb13f8qHuF915nKaUzu65RM1
SyjoQajPzpKtkjuOLLh7nvqo8Xph0dOgPb4SDci5IUfYIwcDsleWCivbKFV3g8lnEwc4HkohUEhY
ig31QVO/XZ5GbgnbjVWgGcAabpeNa92i8m8XXQuTjNmguHH1GbvHKUn62+2R3vp3s1/s3/8ATHp9
rE4Lh6Y+hsBg6uZ9QqWxd1gWiiNXnW0cp8sFBxXROdPSEwK19fO18MgcvZEAF43yAdbwDvGsGMcv
KEChQf6bKq6IOccoA/Y1M8DEDCWrMkwh+daP9ukcBgzkSCjgblAbWfE+Nb1CUI1Ca+XREVAHIp5w
cOZL4QO1poYEQvkQqmvZCLrxr0E35d6W+F67hmgB8azOx14KJSYBgOF29XK4rTK6jBwbdXz2suNF
AIUSJan2avvg4JuZaksjMwiZe7XrsEnmpanc3dfj30DBFWG+1zRgVTx/8atgrb4SfFbbOLHBVbbP
WEf2JEnS9xkQEYDCESV/Dx1FTtIQ6Xv6jqFijAeDo9tnwKWSxTF4lzt6/54FMXKRJutSwtMB+Y5r
Uv6Rr0hUqZp8URQJHVYK8Qya7F7ozLgZlbheOg3GMKBR2giX8ANy/55zmz76d0t0zxJ2BbujKhjR
aRS0jBwVss0rngqnaj4Sp5KKqFj8HC0qT05OEz+Av1WEZiam/l/ZRU4Df/sx4n47P0/5UtfFLdgf
As46Lqnja3ot35ZTLXxwrO5GFaqbYVjEZn0rwq4hFzgT2zuYZEBZ4PFV5bapv1Lw/SN45ulm7MbT
A6Zf/BO7djQ1wwPgA8odVFGmM5hINWAZUYQSzHesdFpRwBTWm8Fm8dcGNxvuIiHGXkLjPKnHVvUy
Uz6e8ibwzTLjEWLO7h+ClRTLJhVSQBk5xaX7SgACqwL7ZIPIxMjpkm5htimhdbBHIZFGZ4QacOqe
J/qOpNSEqE+VOvO8iB0DYxDgsGn9fYJxX4s83YtVLdNCSZ3Kmt5Gt5eucA5rKlJZd/8YjwifGsJA
jUBpQLvo4AX5aElWK0/umVR1d0vMnZ/Rhh4AbTkOH3yCwdaRrIWD/+ztIq1E+QmqLg+/zIMYMRV8
DDQlwMgkxLgyXfyqLkpUoLmVTFUVp0kLOJl7p9Mcc8hG7J40dmd11XOdSGxz6XLcCJ1F5UediBfJ
CPUyCjbcUb52f+i6vMN3uMLtlsHpxffT6KzYEhSaP3BwGI02XRV4gponeaTZXS9tiRxCjD8saJfO
heri9y1cGu+9BIRaSGDg7irxKMOcKUsT4MLsZH7YRv5bEgMcJLQTv37Ta+vrOeiJ8Ii/NE0kiPV5
gNDDVDr1rrCV1vQ7DEtmhPMZHLAtQsOERz9cTZBKzhSXmFGSiB+8AS+D4Hl6oNoCL+cde2s/6xDM
EtDm7SIoE9zXDYcNOQYzA3tqo9CSFZbqw492SQ2+JSXM08xDJJsoj0hojzzqMQACWPUdUpzimQrY
KTo1r91xgbDjjehCD1mZKQFWTC502HUoxgO2ItW9isK0LnLzy79Ztj2t9i4VbAsNecgvdluxYXuI
T5QPRWjaDUFjXyKOpujaAARw6EsrV/agdOf9fqFJRSh8EX/CJ6WKLy1XveBYEehUumoevNLBDM9e
N8Ha4WMG9D0EH9bO9JkQL1I7ExmLDEDl4IluYZCncfumeaUB00ctpUirYwy+uZ02E3qZ/Vk4M91H
SPT+zvD78GS0jcmUYmIt0c+hpo3kcff08Y9iGhj2kUi3yaTtX+VC9Tr7u7dE4AtoriQUVHgNWMSo
G03UkfPSbbm894DgMqXTFnt08ohD2OP+qKScdq8cCd/xkX7qnlwoi1DS6uU8Yt5Gk4aKLH+nD6Cu
K+aNYraFenv+qQ3lJlV5u2kdqyQIpHFiK+lfVJJmRuiLmxXQzrq4z/Qfnq/Zd7q3h2hJrVgqzi+l
1hxOUDOXklLANanl1r4WIf5YhuMgrpn6GUbEtY21ky4C4MBK84l4KInO3K/vHw2/ZWUWSREWhJOc
9OixuNeKpwfLhFyLu/UdGXUTg2hWBmTN6gCOKTKbwSc3ruVttIlOp002ILUE86iWSnaMMTR2/U2N
kciOn6hXTGfz9m9L5FJqTPDg8HwFPBB/9cb3grRHytASWtLclwNwfnCg6gr81BwhjXmR1Wv+i3o2
WDXxrb8Q5mN1GCF9RBQQEO87kaumJPiIyACgilGzGNoFwqdNkjnTwoSFyLlndwlz0gBxrNzam1Rk
Kth+UEVIiTvJwvaJUOqyyzz3tQtfZj5fuh9CHQmS6087JwHBLXPDx7eQLmyp8wTr9tOlxV1SmLvz
ytEMKGsWvzC7q+aC84jcOXsOdDecL8wp2PDPX2aisv0RTGW5R5iVtuS0x2tbMPiNG7fFl/Ky0hfC
NEx18+m3WlVOjlSzc+zDovAh1mxyKB1QoW26q8kO873onwrSLRggGWOwRub4ZIJyHrQhXuDG9bHK
ZLjZmwILqxBZ1uQTtmlgSrX0MXDfqv6oTh2bO1RIXPu9XVsvNnq3xaZogkWh3MKq1ehASlIS7K9G
tb0tcvjg0FJ1C9UhXWXQv/QMbhunnm+F+Xu8swHTNTN+zuL4lnJZLgfpVj2gn9fJf03vZ4wxihOd
vJw8JdgJhXRdXSTTAeqkH39aQqvnZVe+KRVycd7ES5BoLRHLOmFPQny53OjOFR12qXLrVBgdydfX
EXa19vspb0p/irNY6Ci2AHw20UunhnWpG9pMpTI+2og5mVnhsXQqFECJS0oMq2EMmm4Dvz/dOFG6
Ly698iYdTcEsoaTLO/RFk5CqE3F+30bspKbkHlTQhXFthClFBLRw4fb6b52TtxSS0NtgjKeh5kSk
eAA3Bk0DcSeYE0zMfFNnxIMd68iy+SH23TEG7d7DraXQdJVHcFQ98aGMNo1+QzN6a8LFurPz94zM
N2m6+0HZDdZHDOdB6qoaj8pRJg6ZRRRPDasDKbJNbKJgPnUEpzU4W82SvDVz28J/UpRFnww2Y2QD
3RCaszRifpzo++25drCiXQTALI/lBhw2NDHGa6EQow5RwZ3mTRhWU+h04c+dbWWQzmGT10agyMLN
Yqx8MDwx6kcPW+vxPwC05h/5IfNstTDvx5o+AodwrHiRUQXs7f4NM4YbQpM6wdovzqqnXSPgeiIQ
1B9U0yISR5ViXrJre6FBluSL/FYNBhJWTMB62WjKZx0tHYNi1fhc9603P2AyRwgH8IOAeSCb9Ue5
bEQIkOMkSFN85Hd6HQadcj8qhR9ISFXAhc8qT3dMKhoi4vsz6wZCGuNr5WQTWfIt7TCZ1sl1FLP2
MrsbwLsijrsy1UczfQm5Bx9gEbslFiz8pFNc+AkCNCLt4JY7YuvxNyxLI55e9JlUwByWVTIsEppO
BWd3uqLGUfGnra4DK0/RT7XQxus/dQO2xjMH1+mzlZx3RfJDro1s03wI4IcKzBbNgncZl1NrFdmy
VLMJw2GA5LqaTXRvoGXswtSM5aqTYf3vlGOPmnZ7CtK9W6hLC098iZVXBSHefgEhih9WC5L5a1ov
2WnLe3Sq2Q6w6HNjEwcRCAzMrnsvHiv54pfIB6LMpSelgRIfU61iAHbCig9nLCgz8gR2vgHjcIpz
CSSoSPdx+3WHiPI74HcZ5de6U4y5xaHBJ8aMGN6Vm01hJH3nJMqeM863pQLFS7ravJmGT3mvTdPt
iX43rXe2F4yz53sCHrpxBzFCwezzjhCJjZjAKYLWtyEMYLAaqv3RuUJ5aNImTMcBEHu17iK8gXzR
jp1id3u/ayf8VQ8BtL9///1nZmZ4M3rzhJ2b1VoThgMlYQh0Lju9p7odm/0PSeCpz1TH6j9QTcIr
YOlOAPWbJechc4Wi+xqQfZ7UXTqPTqdC5co6gUbqrZI3K9MH6rkqguQmC+FtyBdm+Z02ONn1q7AO
gVxhA2rUlmjCsds20l7rOmDIZmZ7McQEsq2h3e4KBGj/vkUdfdGac5PS0KejfScOgRbk24tYpaXz
Y5UEX6mp1PeVlsHzW4l/RVEPE/XN6dJi0Rr/92DaoCLAmgbFkk+vdoz93AMHK/cGp6wwyphhgMwQ
p3DCaUS4kYcBb2TKjERSYRWzYxrSj7VPrjk5h+yPSG4KV4fh/TKgR8iTfwCqnBScQ02DY0ANBS1x
iZ/JoumgJkUM7YIs+eyxA7bFZrZ+sbN2AzMi4Djbtv1yNhA1Y/FX5PWZl7CIJzJU14fiRiMZNGvQ
wRsWg+XMLpKA/HzHH+nDmBM/34xSTFsGiOmum0A/c6vq/rkBpsNiumTXdBqhfRsV6cp6Ey4uHqRn
QkBNYkCXNMIoEn6SwydlSZ857AJsfY/1re4XAeUkMnmWq4BvrB/cNiqNz+sWemJqXId4s/pFUOUv
/qyKZgO9AwIQ1YvwA/Iz1J9HoPlvlNRtjpDkwcUBOhvKgmgeXKTztsUhd/G8irr373SVENehV2LB
NsXJdjdlEoqot90yssX1ZO9TRUaNdZNbsOBXs/tPBrolQB7gFyTFf6ij7rc93Y8KZvEU5sDMpHfF
aTc98jjBCcqXeiBkZU6WowgF7EpXUa2K147Uxe5QrO8l22AZKthYlNXXVDAt/GUc4FPf3hm8JgQs
tTz/2Wmr1xpHhP8VEGjx9+mArYQZDGy6tKJXoDST0ERrzI2Kjo9ZVjqRYlsADIiLm1chzxlcuAnI
8eCRAjlFeJwA/+T3hL0bjqA88y0WG1hTksgHF4At9AxYtejZnNKTyhBrZ2Z58W6wnWeVyh9RrmiG
G+3JFIOO7L0qxYeisZ9UI/mq6OFcmhXmAwA34hB+7AzJ4WaXuQKq2l1VgrTyhc63RMuZi4Ss0OFM
TGOeOe+y7jQuzWF5dyenOfSJBvt/f1VXJxJ1hvigN0myQAA2ZpljDzoTn46tyRc8K4k7w7gHifXG
QhZCUpC6n2SBS68S1Aoe1gUTdYpAYeI3PCc5Ufw6UuREOdVPd7yV97dTUreqnH/y+YamRRl85j6q
RY5TUhNkPonx3hk9lCMW79taAPAjrH7dNCqwYaeKz48SxqqHGgL8sfZge+ZchR5Fm/TdPPcKYbqS
h/9BQ7nJIctofvbPrCtAZ1iWIrwZa1CeZ7DfyCeTAVM7cal4M3m0LaQIyw0pjKC7cdIDWfm2bvM+
X/BKt8fa1Ch7nqmUPCr7wlQMAD9yKWqAmmKKG2XoN2tDbksoP3hxDmnTsdWoEBt/pFXlHRFmmYZo
bjtMstVgy7JhRb7umL4AOjsgpj7UUc/EwCr3XHJcUz5p44szQJ4Ivn4I4CGiRQyBnZ3FmxwF+aHK
a5JfwZclhs1FUwsJVisuVtm/CImeF77fdzAIGI62c8pinBd6xLplZ5eE0hC0rWI0vTrsrQsNiw25
518rQb0iI5OumSLikmOGlDnd69OzT21RmQ4w//uGsS9s87q/V2MQeFXeMfovXShNpYf+dFk3Sl/J
8lM4NT5W9a0c8/B2thWWRDMZzh9eydSlJgaGvY5sP2hL8j7Ki2yM3HIreMCo4U+DuZXY9X5ZKjvU
7g5w6uAlXafW13KFi2wA/cTMEs+6HzdAGOK2dfjoxmkv3VtojKkV/VDiyRjUQur3E7pFV0aMN1WZ
aAjO03CJSn7hzbsPk9u/pw7szuBNLIO7ANTQpkhWy3GLe4/G6SogHFn+DX8Ni5zjVABHHsB7YZzm
8HZ6ov21VqhAakvOVUn2VHd7C+SRalTwrWGMThjQ7e+0bPNt5KWzKqP9Vp9pGdbeC6nwhNO+5Beo
CDUdyZOA/bF9HEGhtixfSNpZ294y3lCkBhF2L4TaiCnsGawZiKPWaX3t3Hg6dY7p3U3b8isZTZBX
VDi0ZLTC8SF3nfqt3yWlssd7pRYKeN29HcsZ20aXUN3QUL2MW03DcEc1xJ9g6GtBXLn3fkHIeiDz
n9g3ns3TgbYLfv+Chx52ClwxX10d5HGdCof+Ng0KHAOpgqe3G0eDEBL3p1IPPnjE7Kc6t1YE+bee
pP3sokIiTyVC2VJQhM7H29PP+W30pAWp/BySAczHOYtPelNmQpioVw3CzbD+0Myi5quCTPPIq/pI
FycAj6ikLiq7t+AEqB0oKTuRLa4IyebkIsgmiBDBITvjPPEDPS0emavS6SpCVuFydRA1kSO4E2Nx
uUc2fKT6hRXguWXI1OhgD6MaexH7Wqyk4b1mHQb+dlc5BQaUA76i2KCj427LoU54X2oYUbECIf36
FRAKJaIgSz+/vtfCy/mrPCxN5KY8fJ8NY+TkzqNk3wpkpzvjzVA/EcDFY+Bu0k/0aQSlQACfnqdc
FG0wEvHElewRMEy1RtPD2bCf39FWdhUh4pHSc2DSEANXaM1kGV50Bo1126DJAXPRe1d/lKXd2Dx3
gFNMPudImU8xtEHmAJVqFpQAA2LfwMGPwmBMLeF4uNXJqLIukO49wVjFw+8XSEmQSSsDyb0EFJdm
u5w1MVCXx89ecAemV4et2NLsXt36zNZtp9pkIJLPmfnw2Hei+dhLp40Sa9xsYBlnwVS3qzwKdStF
uO70xQOISINde51U+a7bBrydgWX4p/yK3abx/RWeUUwCrpA1Am7alzP6t8OnzYUxPJ/shT6O3Hxo
FXl5bnDqZDBAImjy5VIcrk3uZ0BG9xYmxZGzH6NdDIxOc/xrGBSvN+40nhtixpw83SX0qHhoFDuV
ejRoXv1ikr5hPPG2bFTH5Ct4hHJ42sBTXioToPahhhPeJGyO4ZaFTWf61E1aoV17mZXpUx3t5dCF
mAXdRBq1WvY6n1I/ak7KpcAeOB6U1MRK29qfNOYGfGn0c9zDS21ujwuCyaxfJ61rgAryuXkV6dPv
SUL7qIuYpAanvqfkABoSPTN7d1Mztt0jRMa4LW//R0M3Y0AQVioZBm+V9RJAkj9F961mnvsHgKjI
njcaBfMamg41bY5QqiFCS00JXOih7ATSGHQaeL22SmpQktqiaRvA9dHlusJep2ort6NsH7WngHQG
PF/Cjqsod/PU4l6YmnCPTcys0yXxHy+WFpAzdeZgPswPwx4mwIsrniVZ8FgRI7q+F2r0MWS2VAUK
RsKychrnE/KoxEqYeQX47i2ttKqQCel770OYRZzO/xuQIV2Lz7dPHu6Tvf42zo2GsT/S3BmHXSef
IJTMX8gp4DFZi1hfZPU5oTvKgj4ezXpRTirMV6RisEDO+ACjVzNuzhjnUGCnB9m3aNuYhRv1qtVE
2MFRMdIPT6YSbdhfQlYWJJvmeFfmjDjnuO7PYwarD4uDKBCp0qJqGEhbQZDuOzLXByHDtMxhqFN1
Qu39AqFE23gYQm/iGDvQBAO3IpKgb8HYbp3PNZE9Wkb9Luf5nLLRmThPHzZ15grvXKTguCn+Xi12
5YEUlHcmncqaFNATnP8EagbILczgBo+JkKNyt2uc4wS7utre4w59IYmM9bObQhMLcCPA+UkaU8YI
9DU6ayR061vAP5ybCqpeyQFj6c2JfNOPhijQuSpEhC7MJZ71Agld+uR9/trOct6CNU6Uia/f6lrN
yz2sHqt37ivATmuAY8CYkJOZw+uyrZOxfs06zTDFsJtCHEs2hxaIX6Gc/YSSh6bXGiwgGTdOOSbP
E+noL5z89Gis3sz6LUzqkMG7T204pECfcbpulFSIlg89TsPiM1BDwFdxpLr7kw4VuqVZdBNY06iX
wTb13M18ntjQuPqchd57IUW7RxS3oeVxHJXzHUr6rm3Kv5Qz1CgyZ2bo6dOvQlM/S94mYLaMQjEP
O07zu9YINkM7dGn8SL4pMf2DlxmA5vuo9rxCrL2FPuu108TlcVRIBrLIbHyUGMe/iER0RQ+mh/dp
rE2KEJJx56moHymGvW70iaY7tNZyECj2dt948GJmFhZCz7XMFz9WywOdnGJ42CUiK5l6HPmLhWX3
OfhS0FnN7cUuZI7LAPMX5ywdFHbBzHTHZ/fL5/ASfq8Yf2K19rt++Pmz/X3KagDP++Ctv7PRmJDb
Sq1/mkxcSCGq+mlsTleUVSeC2NRgbPaSHZxqOq/+qUbIuAVDuBCAoCH46U0Fju8L8OXsv1/BQPfU
9f0Vrs+dRiB8THb+58ms1n+mf4x4MzC98ayggD1cUeIjgWhnf/jRyNwGtrZIWJtXDDsIHn5LyRrn
rFmC44bYAPW/OQzRidX24OVFU2k8ksh6zKNtWI7o6fzw5/qpNSG9CKq+WCJv0ZP7D4xb9eHtaEpM
Cnxrdbrub577AEX3d1vdfCozprMsKaso2SCx2OPUcpYEFEwskzTVr1D0KEws13+zCBracwtcngJH
+8rZp1w4wb7wILV3GndNss34VfrxCp8SBBleKK3vO47WcrjErR36GnFkmyog3FJxO3o9F6LgQym6
6BmD1o54dclOX9ZeuiTBJSlEwxK52yVaRI8LvxIzucPNHGo3FQmCDlANFumqkG7x0Z3CGy2OhART
f3IROsru9EHtmTzzbumh6YNUYyEkcTm2AkLxpXjheXsj/9BVGVUf5s3Q7bbR3Inx/Tvo3DNCpyBF
Zpmg815e4Sl3tCP4kSmQh/Doiz6FYvEgEPGUTymZsY16MHFTups9sHv8Tvi/szTf8wKp3a+flrQT
vt+Jso/0cb/Eow4/ieaAPPaDUE7U9NuBbDEaz3N2Ho+SOn/pNgYk5It7smNVg4mgxYitHDniBaVQ
ZIN6zLyV9Rr7Dyc+9IKCDzr2b4zJtR3Gc+cSpcBvEmLSSBPfvhKwBAagmFqfhnKyHX4qutvJHjiO
r+OLJ/JGQLtQnwgRQfF09G0aMrfy1EBYEg0JLliBLTnT2RKdifD2vkGosog4O3memdNut7YZHWto
fEka0pJI6WIlHv3qjZ3l+fYSVPXwK+utVInqTW3lbY6c6syVmBAc1uZIV5sdUCGkXQQMMkoFS8hz
/PZ6tu6NoZtoDa1v5oMPahSlecDwcKaT/TCsjUD4DMZ76jpUa66pyT0q12ci6LnccUBxgIL/wYlc
cO+Eijfbe1c0clLOJVphWPkBpg7c6Z8+/8VhE0X+MqoX8nBiY8j6IUSkZ782xbDXpvr+Adg/R22w
4zNRGOIbtTFWvk3w/TLvEyrv9P89sjxad65PWgBABqDPE+5ZftzdedwbUZpst3UjLQ1fXVJzimxh
ONM2ZTHYofxLUGfDhVLp0rcFvcbQoFvyb9rHrIWNhuvtZAmLPUBppUohCpiVapu54uW22Qr9M1EX
t7kJrmkY6v5Ffl8ZFIstRyx4Vuf7WquV8cA1p7bSnblFMF0x8nPG9+uMCWo/HxY2SBOVSawjL5Nb
kPuPp26a+xedIX/Fc4oF+RhKYz4FOdaslAVDLvoyzOLRQyBCckrG1dxiggqsKfwu728NDiSs00wq
m8gOIDzLzC03J41/IR3JZZALz3acYOGLLHgtCGepqfnLq6Jw24ZbOsh49P9gX8keTqDf8nH48Ta/
qIQW1zDtsjQdFUDVOaCjhGzIZ9G0CmoWTxr8yCWha0ppyuoNXC7alsxLgSjYNEYOpeW6R6bkiuej
pAcnBuWXM+LZAZCa/gHOAkqyJfnjRGcQCWQFDIhh5PYBtnpNqTtk6aecG1x24umvZG1bYsQO+vXn
WX9HFJhoQtnxEmabIk/Py8Txn0khzYge5dCu+Z0W7C/t+O+dsA5gU7cOZUiprvUWPCbzxZPgReXH
eigyDZX9ZxIwPOry+ZMSQqu14mrK5fyJpMzhm04GjNySiObSyuXREKul7ATDxZHnXLV72uw8V+Mr
KVSwKnoa1NifIdQQSbvMgxcuv3rOrl17MWPksW9Zw5YC/6iJuUq6NYNlUxckiTGjWO0TrfFvqK3j
fJZRYnKnFFcYznYmSVhmd2LH69Gw4qfKepIoIcWh8lBJ419ZCI/zmmO3MSoJt1xkvZwMr8oW62DU
Lyx1e4vOEGLCJJdj8RdC/jumopsyu09rYK3hB2P7CVtfCTq3uTTUk3ngO+Vr+jXNYG4cmj05vB5B
RIQULS8ACzogl9KYGabcxScgCsIubEKiMqYcfbMIMYIHRg5iY9C1OSe3dCyUIHA6GNrCGy6HTJGE
N8ZkaVeB8S/nS9gAE7/tbO/qE3B2ARjjAjBjSfbd3Tq12xAaTij3tS1NFiL2ImGs51c0PXipu077
ZHYZmPYoJqNDdl3LyQEh/ACTd97JKtWHXa4g+JTJPtoXeZIehrxRkgBKHTdKcR3i/pHzkrHJoYh5
deJxcyOGIYUCwQeCST1s35fQGoIaU8QvcZCpjrhmcoIU8Y4gRFrYn1E4Mnua/XyhZbVpq4ACTkNJ
RpC8cG04z1dnR+zUG7Kxe3mwIY8Mmvh73/YBNpXNxCkwPSY4TgNGDhS96zcLAvoFBObU1Kj68HoQ
b6r0O9/ax+bHrRXhIfD/J41JVyAO7YaYo3sk1xq1z0yV+fgtNmFBLMdt+egzhN12e+GyS56xNmz2
llnL5L0oYHfifXb2ydtV3gLotXbHpoLoOSK5Ck6ESQAYoKfe6ECqdFY3hDbd709lvjXxLKpD7dae
P3hAp+lAyCurb0JNkZQKSOMWrvcC5W5NrJzmKJPozWVJRVGj5T9UIhdp0vvFXmoUgG3KngqUfYHd
gBkZJg07UnKzpd+V6cnKuOvWl7zPD8r4hDtSIvw8XWJO5N/BsOIRaS89hfLKSkz8Qguky7uhDx/l
Nk+LaUplVmtnA2ULVoo/CMe8fQCleZ6PasRk2S1ll1YcVYYRW1RVM1jT7+lZe1uuRSsU/pQHokDi
tSxYE3ZzvmO4mFEDhOgD+BCedQz9bFLAbOaudDUFRImhMYnCieQRE6s1IChW1xZrGIL2HeMQoB62
o5lC0Im+Xas3EEUAkj2XZYuomG0LT8eKDWzyYyiUyyW7Lxl8XCRV3Fchwy45AvNajIARwPSoTZ+u
5/LG8ng2tLSLxwFy2wSBKN1iuqOBmsVbCY+ZCzWqodPLH91l8TI3rjd6iMnShUFOg6TqJjFwhqtB
OVVR477sakW7Sbov82u2WVeRgihWrzvKxAZ6hUaJgoNppYnqitQzmm6vTi1a1NAiV1lPipJmGO/a
HzXvdfq3N3b8BUDXbRQhKcCuPaM9dcAcAM51VUuJTXQG5gdXz97T4TvGv8BYeW8wySh9lzPd/bY2
V1M0Vx2ViajT8ISd0A3jh1A/6DTKvgNHNjqWfyKJgDl9PGR3sBQbg3F+zgwLPLYbNiYHqB2qxYmb
XC0iwZ1h5aj8qcJczNdKt7g6e9fMMXHn6KS1f/pgXMeQRy2rd1QQ/0Xw9LGd2JCj5YtG93FE9rIo
KaE9EaRKC+y5Zfm5iYL/rn1PymTpg70U5lv9Ewnly3DRG7vEM268NQFu3uG5Lk1gHigq+a+QBZ4e
Ky7Qe5vHfzrk069FEOy5UFlQGN3GYBR7QYZ0cCkEhV6xF5K6Vr0PgN4HWhZ89h9QR2nFS1jkhTel
DfYlDos9Nl1T8lkaEJwdHIhRK6RcchOodMVpE5v98aISWFsSk1i7+Wo7nvep27ly/8kqKIyiTWKQ
1hapifDpisVjpbTDVoPfuXNWdfmqFe4LEjhv96nu61K50K/hYhid36yev0dxZnrbMUmLqIJQZ9xC
XHrMPCGT+I2fIyIDBei9mFi+oxJEuQHMrQpjSXMi73wNxk4N9JuuKTaun1t/mIN9w059ePbwbw5z
rom9+3sXE83ZpASHV/vA0OGnFxRTo7yo6Up8GfK1L/JD7WWYLYuWTA+SOJn0Z7c14qo5DPXSQSvv
9nvFfeVoPbhmwQt2Qx9hVHPlc4xRvTvx9AjBZ/gwtcoznpOK0U7qGfXnG04iTjp91PYaVo9fanV8
LOMjpdwALUNbWrkLiLTY+CaZhomsTivKxKdjkETrFyuGkKlhPaEPRdX7+LoABCxpmBU5QE38JHG3
dujKOQp9yMC1GQeH9Tp2t55X7QYyYrSzQwUTN8p83k8hFlBbbuACcBm3rid1zvM6KKLWYLdUd6wn
g60EyNK8XhQiNDgn16Y8ARTzFzoviuTmJT1iAAqn4mUzyOTzgRLqiucg89n8uhpmk2xAoop/yXCJ
Gn+UIw7tpOYSQ16Spy6dWIKaIgBul2BqbHM+Xl7coboV9D4A9gqoGHshniU7aahy+jne0URNYWeg
q9LwXnRC/Kziy8tIoT2b+fnFI4+FnMdYV2+btKoOKrBQ6/dXTY5s+gg11lXvYzUo8aAZVVTRJsij
aRxDaHodt/iWvq7D4fcbvrmz1hwa0ovnNtW0MFvB/fqVoO9LyzbTnz4QYcceWmP3EdPVSbGKEAoX
fvS2PbjyOFlvfH5TlfNb7cImKF1u3ce1eIJLc85sIIbbQZOEnmV65RonXEeW727wup2Sx3pHfziG
Eoq/jrswva/SvdGHetdD3YmagExNnLVN8Mkn5aicrUp87grpFvePoiSneMQNd/5CHsE3YVCU1064
ezrg1LX2K/e/erN+euxbFNNtFiQFjFeyN17m+VcvfsJtnVDmWyQuDX8hP6CPnBLMmR3IYQlJNpxH
qxVnOlA/7vd8MM51SIeJRL0SidYkL95cmBgcZqviNtljLrDu80rHtolI8uyYQlP9maeVGBEaHPqB
FxfQfpzncVziKuMHf/NOckVpIgWr762ZGk030AXQMliQf1pWR7BTpnMd1R20QnUnajhFtpgR5kih
s6Gt6YVuo6U1IuCmqK8a6fdSwjMz00hTlOXEY5MsVGUkGve9HDGqW2SnLcaHOwS7dangnuvB9FES
B3TEXnKmhSs4efzmm+XVk2juK7yjA6jd4h9y2mkIxQa4ohnTQyDeuJhK8SfPKF1p+KR5M5vbgqrW
m25PigqhcfPRmFqaffb71ApIn/ck6vCJlb2Z431orrvi7odtfwKIlcnUXEQ21cwe8H4JiVt9vptk
ygqOd0DlRqhP5sv6JTh5h7m85QkoEnRV7H7ECBCKxQerBo6QDzyH0kV6ohbm3KC8GgRQc4WbV0Xm
yHOsgg0VB77+DJj0Hae7v85I4pFwbxDjDstXKVkYM7nVzI75ZJnrDjLX4I+WyDq4GMJXWcle8ZDw
u60tUZKkKEJKkx+zliR95k172opHY4RETVNniudQQvKXvLqWeHqAPvLx/92nmDSyw16ybnGJJRoH
4Opg98kIhnf9JK7GDc99MhaM6kfmqkRn7BrfMXKPB4ue3zYTVqWNKyHlpUgKZj3XgWqrKICbqQ2V
Lj1TQqLKcHAJK6Zcc5i0/CJXkI/h+g9iY6elf6x/W8yUvgL3NY0KN+s1wYrqHjM31sgW3S+ah+ti
vb5sinF0WnJ47hoDzED4+IEAW4BaKjQme7yygkOS0cGjkQjo4yGdwa3MzGry+Lo3pGeqdDZl2Lg7
TzbM3Ah4J+67BSTzaolzCrI1T/PjmjgYpLfZHSqNvg3jU37xpIC27B7G7tBxMXVTYEIY2AzC8NrO
ePHHqRppd6CJ/Ie0kT7MwxvjJrHo9pCFeUbRtW9OMRxgEulUgbr0yKXEZnJzWEZyHRHVgFLKHYlf
E3g7yFOKEeRGNzBERUzrx0rJfN56sex3OJ/+HmcRIPz7de+2YNv7xrVWzmvuJTSbuDo7sJ9B1wop
vws+JZxprIBR2vO06+JtF7Kogc+RXNOL8uxRM4TjfPpUj6d3BT7kJStU9KOT2iSyY2jO86S3tmDE
zxwmJm5VuHct8rOu3theHGOUziklQuNZmFoiNHhJdSJvKDRVM46RCGxljHTN1z2o8ZGDvaoWFG1u
kQlKgQQ59xpJBcpTzW12Q7kMsXppu4wfj2i8XLfYXtQciGU+CM0tIibTRljqBr4cJj3vJY1xR+lV
TjfrXjnG5P8/orIpGxUtEO2Ya1xdZMl55DyWuUTTeRFDthwDRrhg8Wio8qd1mhSyOjLVLfon5HQu
NlRME7j4ZsPxAE01MCEm6kXc9rMqTvwZ18Qzf8IVVDPBXJDbSVcOmiR2GTAWtO1TBJaQa2pbNZg3
44Y+jfrCLG5IBagsLU0ehmhfcCLszNCA6MnWsdkUA+S5JMEHpG7bDlodDPDVpod2Jp6+aD6AFgfI
IdgRr5YDY4eCPuvhA0UZnxUvtor5Ogm/5yAdtcLOc44iRYQ5AnO3Dj0p8o/nwZido7XwMC2WniFe
L5TPi0dQAj47zJoDg0WDdP3QETmlGK56qs/1MBRrXU39DGoxerGNLJawkn+WE4/4+mDP2XqV4PNm
kJgl7pePnW663iYFQUgu3rsbGSi8k7jDWRL5jgQYxHRSE0BdWggvrYTzSw8M8fQeFTJGicVHcDSo
Hgn2c16tZz084rODOp8JQG77525JS3QQN8kgXDwkHaScozyMjryqB+nTEJyt3S2R99y2GLHR1ugq
MXZpyWeWtDuC+nVQpMx64vWTdYssN1xgSi/3ZQOf4pvU9SN9vcK4c7A3xrQtedP4J+6TNSNbarC8
nsRZB4UQMLXtlbabzoGZLWBE6+tpDDqGLiqlhTAglmGgSp4P+OagluAaCqHIYlWtzSBRyTrkpeoQ
NpyW+S4StCYYbh4B4+N+f9ZFaoG+ycKxiZcKMTCw2Xa2fX44Lf3MXGe8TlZ/4rc/m9cahmAXyLDS
YzhICnnVBeTkyORyvhIzhEAaO9j5PoJsqs/6wpVmTPWXqc2Iu8bicIj6wQ63A/m/1/U2KdoE3mnU
lalcKmb/7PWIDqdbdXlzYt1R75JRio7oqKwzbqO0Sq4NGeiyYU6sV6li1TK7tx9h2aM2ikO412r5
hDRqkhiyrXwcchbLzVq/0HNeHT0iplNY1r19ykr2+rChv+7YE5k23GeYXQ995J1xD8AbybHYVcZv
vTuBHkGT5uFZ2/E4UTrONXFJ0TKLvgz9NLbRvhm+31/dClbhbPWbKmN1gjfV/T0tE34KdLa6lX4a
w2OydXo0N7ZJfjmwY1M13u6VAe7nzB66LxyPwtyLUZ4APNlroIw/pOPszKJNengQQzVZyKg3A9EN
Oz/ixCsCuIryu/lvapfKu7XKldZjKwXbmoJtOL+oGVqVQmzG7YTwHJ4kx4vttwogtkVi65g24vI6
0Xrc5bkMCYY51LhDOuS4tUl+YhVxlEMlvaN4LhWGZGXqCtd5cVfcGmjwrkqw3jx5zlt2oCssXsqC
ntb/Bzrb82IEdxFHPn/3Fso6R58sdihqpLjSbqEL4pGbyJsEfvkXY6M+ZZX0LXml0lc+ICBmDo6l
s50pgwck9clmyDlxV8YFXPVfrLKOcQxMTH6NWe2xueuXQA4HI1hPyUD/Y7SgtDbPsLgU/mwtTs8A
z+9+BitrpR9DtxPNyTIQSNMYuC0b5fGenFTHprSuc5TxHUTFMMc1qfxFuPDCzMkRLrLbNjY5qDb5
ccb0Y+orqPxtnFLNn2fLbNqyIr17eNvBCWeVTLloULpBtlnk0jf8C+izlqUlUZJL4zjc/KmM8CmB
PHt9vZO4HgG4IvC+2GK1eVjhWOz18NDSZ4O16LGMn10c84FsEwEnV30rI/UPrJPp/ViaRinnjogG
iM0Tdh7bILqmPCop21SuqmJzLZnW8vYK0x4l3aAtDG2nCHH4pUTIg1wS5sVPpeSDFOYNueq+zqdB
wV5QicZlGiZNGpUrAD4BFVs+pg2TKnH/NcGIovmrZ5+zlnFyBhk3CoFenhAT2IBTN0ZMfQ0umvgO
KwrKroRnhVmxYU/NZLxu9qLiE4oXcrVHJnyKmY0CLlbozMI11TY/3MiSbtCNp00ZJdo4ZiMSkig/
ip3lKnlxe9ukyAMlIs4fflrjQiBXJRpw/CRwV3tE9A4MmZDMPz0Zw8WcuQYkP1RAql61uvesb/xz
HYkGnbur62TIdEFptSPeRk9Td3eUKwXH//m7AbQA52s9IozSgo75tdf1qVlnRCkE8s54FvKz20wB
cAlCGAVo4dcB1rzWksO93r9Wb+PrcxRuJjfI4lLMVLFjUCF0yZIDfWH5jV/FmC04hwUDDq/iOh7m
MijCm1CNCXqC+UPr6neDxBaDwermtzlZEoF5PJqxV4EsZ8atCWxf9Y5fHlU5b4lsJp8xRx/tcDsb
pMB79FnGv9qWZ5a0yJcq77FMadQvresGl4c+I2XKkxCh8Tj8dAAXpqvsNrkUzsYQ4JlujoO7Oq4B
/WDIF2eCB58wd9FkH5D+Q3+Z0uXUQ66HewNiYIfpgjAfzWEiXLJt4Gqwqv0ZSJuEbyA5sGKS/+Kd
OUZGykO3ZaMDbu+mfrKtfh7oH2z1TQRCtu2JZ6ju4luz383LajN/hCGk26z8mmftsXR/zW2so5ji
DTMnGFLjTNcBg0/5/T8GXzrkoZjVbq+etelJ6Rmb/zu9FIorNIZyvBtyTnK2/HUxLapSGIVAhcU6
nhlDhF2XkhWaM5TqQUcUOblBRYjUFZfEnSvb1Oj73oaNhXEoHXJ6k7y9G1jtDKqbIGvkNjsmZEY1
+WPxH8LqluvbdezFUxYDTuDdsuvbD8NC1XMBVQg2WXXC6uVyM/iiAXiVTXiZ9Sh9bmx/2l0nh/q4
X3XA9RdeRBDzlHCVFbL+vxPvzwZscjZ537SBryd8S18/i6CR0OnNZP8Qqaie8DLoqD1HH1Cm7Pv5
5S++iLS34wHh9DoUl4MA2m5ZQoVWkgDse62qAkl6ts+8W6d1BfaFuTvdHT3dTv4+EKD8jBFIE7+J
5PfCmBpxihKHfMJFIVmVZ3n15XUA65X2pX1p6B94MhmogmWfLkjGzpyEp+rYdz02rbpYaDuRXNVQ
OXqrwiAIEBVWlZ86jpQj7Z86U+iDqBWi4qnjzBseS3kVUiGB+qykcXIKDCpFrTvXxz4jDq63y/Jf
dwKv5gdsqc8kySrhYa/eABO25AdxYWsy1OWE0GfoQHC6+bIROqPMjzBb1UBbLuCbvAtaF1gfnNH1
7lt0doOUSwaneFTkMS9K6zu+Z4G9HFzbTGmgdHeGAy7V88WTrkOh5y5hTftklODwdxW/u0Scak+H
KihYymUTHGyN3+z9sAIJodfvfwaRsSzO6ZW2Q678pZeLARHCC/3/jg53rGxe26X9QUZHIO9T/Caz
g+NtXueGrzRyMWZit+u5tH6zUzHPEBsCEmI3/cOojn6x3e+MR8TkLhj5koEppnjySlNnWlRp/vIE
vDFNLKGgcXcjMlAPQWr9pEO5+0ZxqFvY1Oze8stTVfMErg3IqO9UL6rHDFVz7iMIrqW0kCTqPL6i
yNAGgw8FR+Yv9vyOjbuTGj0ZAZSnob+cT25OG4mzC5I4cXFIzC9cPtXtK5lWPYisMRIMLoeV3sxO
eHKqDyDoQtnrp6sWgYbtQDo1noritMVQJEyXmgG+KJsYkIzjvHmD9h1CvMSlC0UxD48x3oNfqxNL
++i6sH+g98KINgTZ7xGvu9fnt9+kQg16oPXh4jyi6WiODZRvRyd2RMSBcWHIMvV6E436I4XPFm5F
WCGIrc52GZRtmmMVhKiSaR9UjNOTs1X7TZm8tG3UfiFuzewEVI6hHt0Au4lcg6I7YvBL1IVDXCFE
szJXsG5JHBokt3R+l0xjvFTvboKOsG3zRyPyaFrJvkNY4JBrIVlCbGC0jueUfc+zU5+bmsk27yin
7peMcLDubDGCiFa4aSxWwdxOLPMi/7npKUEuTe8nGrbC1zRybBXNandDWLZQwQKLZHwGiobfAd76
NR8xRc2UsQ/QlJPjg4Hd1La/Pc2YzttiOuoHL3bSwaL22L85mFzEp2nSGI7d41AFqcXsGBSh1Rli
J0elkUR57khwkrOxqjlwq5hdRgkXFbnUp4fJv8v8XP2Vt5M/dppVYxMjh/EEx3PmaJe6KDUHkeiR
c4T4hf7J4uCHypterBrp1xjq1G3PLmbeaa5ngMPUejkeFGj3fYpo+LBczmqqoU0k9M1caHqUzThn
Zf8hiXkjDoxhIGXM3eyaom3H0TbCNJokYA0DOUOsvxkxxaCki3jI0FF/cuG3sgCkPekFaNXnLGIO
WoybebDHO0waLvrNAWJPuiRaARfTxJrFQa558MGumvaQyFadl0LuqD614/R/XcBdWggm2qQb+BQQ
uUM9kODTgQo37VaDs2wmmM4OxL0VXckrS9XcWY41KkJODZJhmwkfl/Pf2pq6iPnwdLMFXLzhfyz/
tLHzmPUv2nps9MyEZjKe8nKZe2BfZUsGXFAz123GDOOGhVhq0+HzWqsFG2YMr/XlQatYbIyFMpoX
yaUpZpyQuRQjKJXkkP8TGMzlZyOoU/I77p0bMTqAT9ZOcLzWrg+zg9Z6l9JgMlqTXJwYAxaABGHV
1bb0meQY4oJ9SoKkH4cptRcdnrM3qRolW7HNF3/jX8wIsB834BqSoJfGEjD1cLssvWpcdIT26hxe
Vqfj+5AqpTzLawQD70rpHXRALqXycz0cqMhIMxNtO0nR1i8ozYg0srr+RFQD0lriXgJGFknulhKz
TVqB
`pragma protect end_protected
