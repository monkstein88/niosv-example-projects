// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
eWpA7zFE14wW7q+rBuFR3/+417i0lWJAI/uuLYdx/f/G1WagDA7WJzYkGuUbv4VSyMg4UqNh/yre
bV2/ax+hg51/8INH9C3TJFFFk5n9Rc9vbrU3KvdsSmvyYsbXVyIFYOOZNB+tvuvfSgwc9ouATTlk
EmqRr2s7eZSy2xyCmB/wo5JbiWagFw1e/FQfvCHKQxvzxCoOCMsLKXKbqbXrqrRZX32/zE6Bb+mI
M2VyDbFm8v2pBRVRuwCHsffIE+xjKaK7ZdE1S4qpkpfQ4tPeqXAGlGwEzvgBFtoQO4SskG9pleZd
xmx0iIHqh1yIOv9ekx+VCx4bn9hTcwlSIEX/tg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 39136)
GyfmE0l9cT1wAFLoIMBFFjNOeV6Fd2EXREkN5DrdrF3qaJVRXRVjNXBB5W6Fdv34WdJlfJmc7dwo
TxCrfXa77pQkySSWqwt+n7GT9VNhQE+xANCUPPoZOK24wtT8Mu49/uFa9yPlOxNHgJrhQakDobdH
u1aTGkNL1EZec5m2P/1Fp2CQs8RHzYfSC5w1pGXYxBueFLPEqXNWK+okwvL8KpeDJcn3/HqdxSuv
je2o4VdURrA+KkdwdfbAJsBJ82r9g59J/kA9xSMWpk7tuGdVd9R2zKgac8fpAW6GAOOVAW+Eep9B
Xw2R9T+5XGewRT26wB8EBsRgs01wXZHHM5aBbgusZLeB5XNem/Hq7jyR69HZMzc0HMJckMrZ0Ql7
K7QewWTolAnAvKeHwelgN+JZ60SkQOH6eXhs/GXGT6Ht2rResM2MB91AMMTmNzL95pofq0IOhISt
Jnfsi3t5ss30IOwyFPID2w/gXPj/PrJsXc5+OX7eSGTSpdQLywySTz2N73Y5qhFf24SCLPYKxZNr
rIDQqmzC9Q9X3JAVH+k7dYp9ySuvgGLVzvT9h+2vKhuSw478UXDvaTglduaWvpAbnh8TgGu+tiBY
FWkIyqlcCM9CKCth6g07kEMXVFvHXR/Re2p8H1DKWvEWTEge5BG9x0MavDioc2zYy7gg6mlnD8Y8
aCS5709Mm7Ab7yCHUiEzJCP96+BuXEheTSyJmwbiDLkhHlYHyac7b+D9XhV/Vftx/6wvLBGLK/kT
P1LxI7iUln3kCPxPvpFHpJ8VvyijSP+eibQMeG2iTwXi+RxEI4gD8xlXagyyvuC88MGqTBGQGAo/
DnrIwH8Av3GvDLRVFaZK77pqocB6bDt53s9Aj+SWjc3MF+w9rnKIZOv9rDZzUzcodm8sn1BGwvPM
nqY9byaFVgUB8kS2giJMTXecCpbg1y+yO4NtEqc+7el0RhQpeciZo1SgKoN2DGE8o0fpuxsykPua
mliDoBH/G8LiayOEhHeJQWkF55t5YYdE0EwMWSq+YIY+s6fqb504CW7kZlFOuMM0Xiou6M7FT+fk
kjwuT6NLqvPVBA8R42oTJkLe6hD0INv4vsv8DTv6DaEdMgbjD03M1fRvmU5bXDFvrXGWGZowx0Zr
qqJYdd3soo+Eutvm2VcEaEkqECvu4kWbxWEgxQTFC6J6cg5M9g+XK3gqrmdTDswlOgGM1vyESaQE
T8dSeNylscp3cQ/S5fKxtmAtD3RRxTAGWs8fiWx9UTqfym2a+fZYjE27FfJtRFSaYZOLvEmcRwoI
LV6lHsV8Vx7Mi6UqYoLMBZfyOQz7VDkFx80qioqYuI1ZdGtQ9UStpAgjUavNi3MuQSTpNrVG6Cby
Ywa955UgDa8Owojvhy80+YGYZdp6Nojd0ISUd3c7ZJYN6lGJdx+o0M1SQdhPd1Bcx2Zv8Uwq90sV
xmAx2uAiD0hHfu3bM1GB0Plwxhq/WPDa+QcTQ3PryPPqZYrlZ0B6WIIECk+bewyr/j05PDm5k/+E
2oXh83Ty/kINaEUAHdiVSvY14nBe9cq6eZzGTDvDG0gGnbLxMBeIdS4pmOmlBIyHnDRZVNrvyuq0
ZQFwe65AxcIyGoqU2wRx23+70Hlbww1w7H8bO9nRuqJxus/AXU6iV33d91uiXkP94tNT60yUdznO
FB3Yy3Gn78MBdydhatZ92wNTXZTmJ0CGkhRYrl720B6+xr/U+ZsqfxyuT58CPDUHXElb0zzI+Coa
euMFqPKCjRTOw+1sc/0M2HmXcE0qcLfZv1UcFepoaWlsKhhU1TOq57/k1a0li+3dLSUgCKJvTbmS
FwQyLBGHG0XeEf1N9aFaoBbO7VqEWkaiqH/ojIFxfOYC864JTE4cuLXckGGgWPtQGPMnK3CYGjec
FkTSIG+w8LAWBThLkJUrCk254q7sgwohV4w1xu1i+mfJDr0Gqa4cEbToCt20DBnG5MelaI8F0uxp
uAsjCRnwOMObht87egOsEspM/JZ5voCqOXM22XC+gLs+JxWAEFfM+wcO/JIKzhRimQj/8u37sbaa
yGyANDTrORfV4tLoRbmDRU6lGHBCerZNz5lbhElDuI3elHGrFTdLD4Pnd6KdZK8pagUERd995AIS
S6PBJkO0wDGbWsMSTw60BdcvYB2Xc1AVteYV5lYVlZPjDlJYPqsqBh2hAb4Unmuw3eaz0lf6DCXU
74LJ0WDH4JK0dTW7bCzyuAJmH1DEQAKjlc0LMBe5sRmuCnBunvExPMpzp/xX+vr9TeqjoFBncYKx
dEhEQ2bHz1u7/F8LsKKbcaPFMRXlK/cM52IrtUsGdBcGjnbYjh4uyOPoIH52YGuLVEFpjE/s5ZLy
5s5lsk8Y6v7EaiCeldDF9s5y8J7N6IbsMs/pWc1MoP/VkUtG0FUdqPe9h/cgcq0fw+QDn040SL/O
Vpcf/uILWBYT8R1czGxyvwrQF+vEXsbgKshl1nhLVlgtWKDPZvNiUcAoPcrSbfKmcOf2YX+DCF59
zaJtcJoARqIH4HmLRlfKzhG1AIrHAzMMlIon8/TNxI2dxma+6kpSzA2Hh8eXDBpoAysLb1+Q77sX
cqEPsUUxKdz1FTEzVuo6/aQLCLX9Y68naPn3WQ8k+xMu4sPH7ycSWVoVAKnynqAMiAISNTOYzMPv
cnC34NWyA4qSqgUoUyDtTpiYIq3AU0V8tWsRq3eSCJwtBYmZVry4E6Bs/3vRbjXf110LC/e36qQ0
lV0WUX1VKmdE/i7W1y+BKmW4GsymL6pk+hwcSmKCBRA89oMXqZentI1IZTCdJ5gDl61ToyuNM2t4
JzGnVNaFJIHlgcTGbtnht6tDpEdcqIpXg7wDvth8VVeNMNlcvFzSpUQ3d/3VpyWLIvKv9laLDdGc
Uusb7+V9ttaVL0pPO0bzTmQu33z6HSvfTLw9oK50I2IQza/KgdJQ9AiqzrL/yrgTL70fiVQzsvoE
uX/QPJ6FiLeFf6nMnkL6uACMa1r4xqsA+7AWfidEBn94v99p/GXFimmDi1VJcvlCZOvhVVaNcMGI
NPJVLIHUPL1KsKdpg51yQNMr3flU9GsdODxrEkP9GQLt5iAiKXGfM3i0zCWpMBndtUOtFrxF7LxW
p16vRpT3E1e1OalpF82+/2KVBcr63BUdSXhGjyvvj+++kfpVEtTE8BFgyJRs7B15saA9jAyklJgd
ajNpNhbanZ5/65OLP1KwHE3rDMxLRlFWhxO9wu5lMSy9Hthk44Ek6kpIGmY9rl8X5lbmw75OtsnK
nloJME331lLNdwpy3m/QlirNXySRyS3tRnPz3ATg9WVy5IOy1OezhiPYRlL/wVRBeJrIPG1r/iht
uaAamruzkj90zsW8CGRRVYRSUPPsAnDmTigyrbWTAASaTgbHkGceAPOyu6O+QnyBEcRLMqoaPZ2p
73odLL3JsMtpGaC6SdHjSyHG2nKaCHrpP8/FOIZQtV8cFcrSaBT7TLZv4pi6Wp+cxseB3BlShro/
Z9lQKzC9AVi3fZAJQNVjlQbxptEuVu73QRZb001nyAZ3LY7uo3rpq5DrCDue5oYb3/46vK9P9hlz
RwALmrJJO81ywg2mxJrbLwE9utf7dapn/jmUNK3Ry1ubmv6IUcu3tFvA2hVXaHT53HqM8kDObWYo
ZutMvRhJFiFLLBwCqw6GMhEC3ub1vgomv0p8r7YpI6iuwa4mpvbiiBlKGxhiGtaBSN8gXC0ebdGk
9Mck9P+kY4WSbKs5ja5iu5ZKDyM7+i3fJAXjQhzsWPTRoOkgUO/9arCOa2urRTri+JxznxRib6De
Ecjhdm5aQquQ5SMRki2sp3GUFViTHYK0zxNAWSvCAsc7G5sKnsrhRDkzGGjpd+eEtUgBgWCuwN7z
O7pB1VX6azOUjC/AoMSQZa5Vqq/Weo2QLyZPaCbP2nQ8yEjaOabXaLoM0S61R8y/KtHQk2ZyQe2Y
Ivzd/wiKO1Pxk94NJ7p3sn7GPrMsgvGaWsDribr22GUIPUZJEJiOvsPSf4hIZHwEpxDZPdZKA2Cc
lgdHLut8925d8eF9yXUdTK2DK9+sMBqieg12fVIp5CHl14TrtW85v8Wi6kcOu1shtmKjeMlY7iyG
kHR0xAxq7gvJi91Zsf0zqZ2BAm4EnDz971xN4KMQxleSSLKt6NtFc60gmdVqgQtZRtx2myXpJb/i
5j9pMvN3s8vX6siCOYgwlKA28QGrsHgMuag0TqvVnVySSWRpMxWYnxXdh8+lYTXOapV//ODDoGj1
eM0mmkiF8PoMyLaXJvo+BX9ueCCM2u+rInl02kTplgUrhBScqslm2K4v963nZCH+d68i0y03hsGa
09g6FpvG8nZoDTJImkpai8cwXQke5ezTqGpCOXfgftxiD8B34GxLxq+zJwk9oyXkDAZWnOJb0gK7
IymppAebJz6ZS7Z40pYQMPlvp+M5K7bfHkcqD5o7XBSX+G+BeOkwkRF1jAAOmXUVX8YM2RfUMG+e
x6ClDqudqou0xB8KjrMyzAI1YvmXlnhF70x2fx2v9e41U4TQHwJ0gQj1nphkd5DAwNi3b5WAotV5
3Np2a+Q5fFqyOQDhUs4B/K+c6bZxzexTQe91QHNpdLDkFErBmKnzwJEyjQbr08fJsfTrjERUTarG
aaHdtCyHagKK7jUNsufteLcTiqNjqbBpDyRhEhBpx6po8KD/T2U/Zu3C+JifNj+6gxOrZv8a9XGH
FU+3NJ9cABMLmfHlGG7ScD+6JhdxeEloPG+WFsIxYmF4BUbz/q37tt9Ry+75zUF0aiIYmvfXRidM
/OBqI/fNa6jucR8uZfXsWikWNLDBYxscTXuaq6fYE5AivY5iJ+8pi5sFPfDMvJLz3gVj1I7nAFXS
DWtR3Fk1r8ODO3EqACBR1cfvSW1U5CqUOBb5ZiBOvjo/pKB9dl/xE3k0wGmuVjh3CXCUhXcI+dH6
s+hoOHajkq8Jl9kLm8dAgXdOBc3sIcmPX0GiO1+WUdLXEWfaHwcmK8kxwsLvqiYex+alSzoZM5c4
eLhmPezE4CDtlCUZtNoJx+0CPyIDioTyvySrAbRpiPk6xYA2HQUI6Z7owJABWuq8kaHaySmB8w8J
7OVckIn3Nnz3xi9Mvz36TrsqCYQQsYW6zflggDKG1lwhWAwA+pTfkus1x4+6XAI0lnryz4B4MmK5
3TqMGmrpzMJd+KpEBs7JRKWgu/xNGMTWgLnjzaGKbpgGslKHHgrn4mfXp9SAv+sGa3m6RF2EkSpK
9XRlI1fgbTyMtvqk6df+aNrtXelv2giGnl7ONgcW6nYADWT0/m8fZZ408LPAo9RfvbBWncgh6yLM
K9wy1taqgPipXv4MtEWsLNBcOj1h6IiKHbPbkIObeAKa9XONEuCmf9PUygqvxxiRYJobqzCThEwM
H8raI1im3eDJ3HpP2RfdGuHed/SqUJYTlJsD0FAO+qNFmpVKCqEXw2NuHCAePcypVIbeV3K4/m2H
+e1zrQyEnKI17xwAdtOU6qqLXCUU8aWN7qrbT9U6v8E0YN5eKVvHphw0R6iKFOXfbX63L2pTnoD5
ZeYIP4KiN8sVU+6pK44LL5t+FLtKXd4EhoMRqzoEM+MyWpBqV390yKK9Leck2L3xDnwI6hcw3Tqq
Q7PZPTdnPefyBoODwQf/eOCYieCn3reFd+g8GjlBAKGlfLvS5Okz/LtYmMfjVOprHz6/UvOmlPTB
CtKE0LBhmgiOxHWf0Pg3Bzcq2J7fXAB6K07OpMc5W7IZqTJeZhRdc71qE4PNsxrWdKlF37b6QA+Q
b3etbMSUDhQxuXkQEND8W8cQDHU7QcQd8aE3B0qD73dBszgu15lnLBxnBQjCFB0LPK/9zQqEE0q8
6jUw8OhssIZIK+KDUpIrDs4707QgSDEhM7950IO+IDMdUk3yFWe0xyK9DGxJWACsKdENYbxB8a82
DauB5q9yC1my7hO2BMJxZ8b/JrDzEZtPTvk+cvuxjtypNK3L4XToyu78GiLLuPAqnVwPJNK9RDHK
TO1QWNAomqqOJ0RRj32/PCAny21VbUtNnVlCq19vvMnDdbQ3QUp8tID8N9z9WiP0poRrgcxKockK
1edxyZPOTYDcobDtSAPltl4OnHD0LclRc4Rmu5s0uy5UyeIEfURpoaR39ICqsDcF80bC+zkkY+3r
uAX5fCiMxtdWaWtuD7/YmQmiByunUYbgXzcy+CLuIF2EBKjSpzXuGNSSaa3K0sbQPPVOSQnBsMDr
YW1rYt2T7W3HCyIe2wx20Uy2etMsFczioP60fIKDqymsWy2kvpKxh0553MgvzN1olOLopYJj0Tfd
t4Ur0wALXyt8IMWIiIeTY8RfUiC5QQaXLHBfV09xR6zIEDolkWv9CfVuNY6F4ZHyadVAEenbY6PH
bSSmlWVnC8swuU+gjVG7Pf3nQhScxqT93BSucPooWlaPu58gNI5xYfI/koGnF2IfOv3/7crwYqNM
22p4fuyD5hd2NaBnOq+n6pg44j57lF1kKBd+ub9rZNzH0/erNUIeGnMwJP10O4R41S02O1wx0zQj
6C2ii8LNzfTSzYdv7o5nGpVoMQPwwn/IiarGs0xwyh5JaqSiXzdu9uZFVzz9Yl2JlmAuzEANiVFM
QLr5DMZlwTN5WUMRhRd70nuKezohvdlWizOpulFgb+f5CLDyPQ+Pu5UIxbNb0n1si4rkPv5Wqorq
xfNVf47iLSUE0arGFGE9/qKJCGw7pjG4WJ+yc4w5Ex4oYIwHIfXjS0T+3BFg7ikiwCF53M+ly5qh
XAWrLVOvetUgZI3yyfnhX5HPRliZ8pFvD7IXaJkCqovAm8gkDabrPtr7bFY1jFjgiGvhZmjkn9G3
nxN7wdx2t1fy+hp1lDPuuVkyIkwKCkCBdVo0WVlGm9+R9MkqIkLvNAr0SO9nd4wNsjpu27uiV4Lo
xKI435MJvWCKk1OT+YjzWMPlIqrJFcqk8fVKrJf6gRHLWKtrEFAaUHHvivm8Hjft8AZ3V/WLoE9K
YHvIf+InpHVOT+wnvDJiU6sK7QsA9Bco7+hBJhqrE10o1n/cnKiWCOqX/znf0oHzVsrQBasnKOgq
Pg30k0p0na4wTx4eLNq3oxgpOfcU0pxbghghen1+1ItvWYXuHXeKu21aqXxhoMXsjR6WO2GnZGuA
u/EhChxyw5yXDOiEyyLpm7wylKRE7d0SPXNh4igW4ojnHB3qFYIq/U37FpfLhJ2i2tg4Uye7qeGQ
igQdGDhnq10Egt9zJxyc7qvPgdnj+g8/uloDYAANn5sPCbpVQInoDIJkE2WBCvqNbU0hMxvvr4c6
9ADl0yXpMbOQjPnbL6uAc0zQCdR2Trnx3MUJHjx1WXtY4x6907cfKFkcLSNpGVzK+LNHiZoUpHh1
6WB9xYXNCSmNk5hlhQ2hq00mCevgJxR+48LSE2fxy3Rzwpt55e0b02nCIMi6BnEykdM4RVGA4foq
5Fk8NSYtADHS2Uu2P+YklwCChRDssjOgAgagnlo8xNE5p9uKlMmFMd1cfCi96Tp40xoGOoppkEaX
r9SB+egODzXC84goLUK+NaK+s/uZy/oxdn6y4Kz3VmVsSTBbyX1OW01LYNeJb7cTingHur2wm3/x
1TzNYh9likuAHax1Fv2qI+qI/e03cki1BtzTx8wq4MYFdHwvKJfBrCpWh/ssdA+KOPsuSS+tkPDP
6FKl2Fqsvc4vWDz0+A2e3TXWFCgSzPjS0579A0lsENGy97RqNphHzQcTpdIvBKTPIgI9fNZrFMkE
xeYPcTcTeSN/5Ry0lxGHQAPvPkopA5lXL1PviPE0V81DA+Wrbs/Gy4Xc2ynOjBZ6eGGC/JkCEiAl
l+qvTokBgjWHWNDR5miGB0Jvu0BBKjeTo+PES3rJZyBYTszvC/LDnANLS3EJE+SLBmbB1aibA1wC
ynwRnKaOusq2HgbnxMqQ+Di3CSSEuxyLasTVN7at5wwgLrnp3oOI7+VX+/r4EuFqkZSrQ+G33966
3137Oa88HuomOu4Dk9/jYF6jA72VM3n65iFBcRzq5S6i/1MNfcogrURtq7tbUmLhjL7wq4xTQynP
4G68v1F9ADHxKmk/cwvmdtlEQjoI4Cutft8GptzwASACWUOLXMXPAG+XEAquipuSucdawVfkOlX+
tzfoB1p3liqiOTBxeukxDHxcNI7fJAmYLfc+eVQ8KKq+rS6W3goQxQ9mgm/1w+0Dm90khu5ZCoLp
CBJchJ5StbggQOlxXxOq3euQo6RcL2g3yhyW25EXpuGu+C8+SxlqxJnmO7ta0kxUmx9+na+vUiA8
GNrmuL6ouMTmd1v86WTzGtur8j61SJPDShSdGN1aJQr6GZXTO9/pW4x/hEpzA04pGj7pmLe0MSjb
ITFYyANJys4oc+rH4InBevf45HODH3CYKfy6TDhE606zY/4aWY8hIkqQ6Oc8dHyotfPys1QZG1Eq
AfjEwOGpgHwm/ouJ0+RghoHtcK/ZSP6ADfCh6YpJcAhapcJqtw6mtzBVUPkJs1p7mqH6zw+Gn1KH
3+NerRQU05+LQlr7IZfRO1qPHKOcMp27ibigwfft2xROCXJlVsO1neQFmbVuJxPYVw6dqVgwLTJ+
P9UBxZfmSwGBTL0ZWqEEB0BZFOmrz9KTJwDbWDzZ1Ms9qDehR81VJ+YOArr9WYnoHm683Mhd6aJm
LYQwiZ4WCICqiVjViBfFnnoaT2G+DpbcKY5rUrNMif8Fh+PIuBU8NyhnhXAiLWKhPK4E76J/cV81
JXd1YG17+LDo/ucIgd+cELK0lFZwPVPw7WOtqToL+iIh8eRloRKyvNs+aaie4IngYyVfQYywlMvx
Kzynd8J3GF2rOzpn6ZhmNbRaVoqFOCLnxrfDo5wnOhOq3RPkysMIIy0dtZNEafJSRCxZy6wpbzYS
zl0n/8K+Cy1iuF4EoTCCgrahTOJ93hvvamh/DIrlcm4vY5mV60w1iFIux0o83WfbYRUGi4p51EaG
9zSP5sZZf1qoubt7oCd/URLMC0zgZXroXbTUoZMZkT0B/LCg38G10HlKme5AJpiNn3aOapbU5WlI
jaPHJbpGkDmlhfCCde9PG6hIsQp3jhtBFaPwqy6ExZeI9GpSX7wHsZvqXA2+jjcL3KD1fwPXQ0Oq
wljKBEgYAxxglJ4rfF/wzZvEw9RAJ1UM6V00R/TmftN61auLziNFve1kJdU7V4Oyb4a5v0fcCkWZ
7/YJeHen10qyUlrZGCnIAXmQ3qDV6W6YDU/T7n8aJo2MDij4o1b/yx4GyeJlWTCqgPKxFLQFWjNc
aK7Nqifmw14TDr9B8iJWBFqxJZZ4OrxCCup+20PdkaPZ+qI42Ms3R59n3eULGp2QFYdZ/Lt+x9xd
39Hy36VOVvhnsft326YwcTr4Eakussq3C7kaEm+ObPJmqEni3ua6hD5Keb4Ux9CwaXLKJvmOAo0+
h1Ue4uMkKy1w6m7sXCDeSKEUx8NcyWiZ1pDslov/9BNMfK9/WpNyfaQdr53DfOiO6mQircg1L8p8
srMqS0gSFHh4kubrw5KBBKzmJdEB1WplUz8x7AMa8mDcgxALetbAAC60wjEnYJt+BbnpuNGtw5ln
jAcO5C3YLZyO2B9LOpH9ZFcbAMD0M/tTZQ2dl3aJdsiP601dPHP4/5m26hSa9tRkOgc93cIBk/O+
DOee34KSIVykoyfnDu7quN7gtksaETdhBbzyZHchGWLW+y0Mbdjs0exiPhIspN4t8rcpzp5zz10c
L6t5sDrSBAjZyjwnJKwi9mW3Z+R6bJhFDsVoknwQc0qfYxysYruPDRc5QG25yOQZ2fldJvjJzSIE
Gpp7YT14u5UvS1xuOYSbbd9zmJthyGbzHOWRdtpiYIFHXjfDNZRJtziHVynEOGYWTqB/JNO8DoL1
8P8Ze4ZqfNZy0OOomWMz5adHEGi4pO6lP2foKNni+6Z5zSg1dDrwZDGbnY0THIY3OSPT4nQ4LWLF
Dy600VYyjZURzw3ALad2C2oikZSpk4doeo2Yx+fcBbD2uvnxL9xuhNps//K7Duz63T3dJiQw0+Ef
yjqb60Y7vYwVc/eZJ8fMeuJpW3t/SYABj2jRFwhlfxOSVPG11HYJss5o1g1GLHBhW7f9nsFVYIO8
76bxCvCGJcsJcSbP3FtEoYtSrtjpBtjcaGpUxYUZtsonqYM8+FczCS8TvGDAympisod7xBVgogdT
Lt6ops8cZ4EBFA/E0jh3VBU+8vkSkEUCU9pfwezCdahPvKfjQ1IPU/vGXLXnky+7iSirNfj489OE
IDdqDXLer289PPBj0ohcUUAow6HSpJNucA6u4sEOTqsSh0atT0fNx37X9/99II+hF6mQ15tvJ6Hu
EgDdhID748v4tuTAVZB6I4EIRqy7SMXk3hghliGBtXtDA+mjAJha96u66S/U2lh+8og2pBbooWRo
dQ+1wHuFoSHTZlJhRFL9+GLRZs0yM8JdMVZ3qQp4t5u+6+X5bUWUNftaHqC0pgvafBkU7shPMj5I
i3B2bnkIHo2N+CHOGk4QLI7eAW/2et/Vy5QtuoXGS2ZT6wnTXxgzYmdTTcL464gTrhBPtUQW4iYX
lOOwcfc33Qbq6j9Z2xja5dG97ahjBMWhpnvLj8VHxmPa2u0xgq3fE3Mh+Mu1DAt3/wX4VAXQwi6u
yPV3xoWAh3na1A3oLsXkVdpe+KCpb3ecFcRKyfgASHJvnLD/itlnrq3/gzumQjv9hEAsmIh4PIQr
pftzd3wukBc/zsfzhlMZd8Qq3W9HtaxKtolfWg1HcjVY9RTrPsM2Liy0PRbZzr1dMZu1XLT8SUiK
rw7jhZrWd8VKL/jTCd819rvz2jeNioFIZ60k/JV6BA/UzxXuoQABI6KLAdMDYZYYPuE2uZnd7Miz
zaR16oBy6LjH7varFvvyWVgObA0m2IzN0vKx1M56S9/JF5JWQsZbiwhtHtMd4h8hg0G85Hqbyazf
56VQACOobJAWjP4kGoWQXyyS+b4WkPHpP/7yKZC4WCRwP3ShgCuI5Ani2r7ouDVraLJ8UCugHPEV
dJB95AUa7XuNQ1L/e2mfd2Amy1Hb3JY1VruUOFkMiQeL9dDP66e4lx9/uhs664Ggva09zsAi8Hb8
uQgwBLzw/lKHMonqcQr7SIJ2uyXANldQUqqk0YXWfUMgxgKZ+1qeV3kaoHD8UoeQLwLIJEkjt70e
vF80Qjl6yID0Y2gkrYP+cg4bEonAu+l2GUsbNiapaz1zjYsaitRTkX5nne7V94ZB6NFbrwVZHeQP
LhOjJpIo691WbLiagQFrODKWDZL+FW5ujWEuo4dTw2gkhucyQB2zc9QIDv6Hp4DyG+XdiM4/+oXt
ANY4a+blzKNErdM90dUylNYxKIYNs3MaqIAPLH0bxsAVTZyPOuaZIGnfN98qjNjCbTlMpUeo4hmA
ufSDs5I16xhbN0Y7MUq3wBpIs9AvQ17HPjm1UA36cI3Bwt1TZBT0ebcwCOh+8LiwCnpr1hgn9Kqh
iMNCDlt81aHnRS1bGdqrLakBczZmp2zR7M8ymFwRx5mV7ugshxqfh68iNq+P2uuQry4pj81X4tOs
VcFrvN2wq4WBjR6YxJ/fWGyB2xPAuOpufe4gWLm/9cFZC4nvT0OMDsVE3lm7LNRsXPDbJMCn5Yha
16ycZuO71bJ6gBRKLEcXoU7tgXCSCDAoYVR4phcBnWvudDYnHUEapw25KxdQjIF1vuEFFFdfpWKq
58rAhUN5Ps7kWyaQpDGz2tE9+U8FjyaJKjCL64kWtcIFEO98NQqUxDSK74Zt0pUntKN8xJlCznDr
yqB+uqj/E4dnsjazDK4InmxXL/BWzUeTjQMHnKyB2/AlJAJ+JY85Z3FBHBUlSWPheb8JiI8HEnlH
Kta5cWNEGGDdYDomH4ykWmp1j84pDz1+iVeFjmm1dDlD24z+U3oAosN6NDIOKNerMIu7XEln7RFt
hW52ZeRK3A/nm6u5mNjeQfLM4tShlhW93A2G43xbAC/fdvYxZoQ/xR9UPj7OMB2ys5QiumYQ8FxR
P4KDg8IBfYJXFib9U5OnJIdojDDzWCzaHxHEoDtnWZRhovk8fqPiRJbZAlXI9qCF4R0GcOpUFddC
67ucqjR+94Qm49aHfMwqJ8P91HQzNf22+0XvOLoeK8aR84t4SMm9Hz4cmo0FoaG+cb8/hba/Byiw
gIp06JCE+A2R0lLDeoLM/rPxdxYpTQekdsl+t4wiepiHbYmXSYts+r+tVPkCAh2mcxzv98MxJX2L
7eEpGyFI4aYeI09VMS2CZ2PIrhjoz/Vr/4MnVaQjAQzigry/J0TmyzPoszB/1nwU3/87K2cVtJt+
FrP6daVBQKycVvKUAOd6p0Jl0pxNkkQNz9Noq1g5rIyupdaE4J6hZ1hztF0Sop3HWpMAKNUah2Ca
EZb7ETfv/je87U24KA+MrF7cVYNN0zRI/HY5hU4JiUMcca/8Qc6mVgYqWBG/cYRAnOPOqKyU7tRB
+G1mc9RCM9AeKMrCC+n4hFbPVUcuAafh5x3pMl21AI4hNN4b/lal4X/SO+qVAuFRwu18c5a7oFWD
2q+RpxQ8Tvs6aM/qDsvxE375sCm8wqVlLUko/d5sdPT9TnE7X3i4F7j/zJ59j+KwLUJrUqEawONA
Sd4f0lOtzuKDvz8J/0vPQgTRFh6sQC6o3MOKdCe9D7rLyzE87sxHX+CT3InPB28RUSJ6WuZYqCW9
02PJE0AaV9gjQ77T/5o7W9uDPXvRobMmh/o/DCNz3+rPDGN6ScsmDtEJ3N41esr6CSGtLLnQO1ts
3g4PkHCsRKkoN6Jkl/28c+j5rx447+6UNK0yIj6NgfzkpdDwN8cb1aZ2RjD1mpObNBoqwCgwMoZk
kUpr53YfXnamYkNKaYUtAG8dR9IJjxKeWc+1xWOCuAtTnup+4Kv2Ls6zT9y5lTd9AcyhqqW5p2dk
00YWr2IrIjAp7kn6w3cSwGUrcI7/ebsKeOjjKX/nYmQAjlytCwzwRy36A6VgqUHg1pDo5UOyK7GB
xn0KPTV8oQuJ4h03WLPCQ1gIuqtOyaVsreDlNesIlUDfzaw3I1fMx9zBmiz5clgH3jRbzgoPYRSG
0bW5x0mUlWzOh8oGbcSva4atKmBpNr++CxMwXh6704oISTGDdWANTq0TneZinqiUSW7FZT439KUs
xjp01Rcb/R9GsxqGgJFaCUDamWNy2sKs3LByamHxTABB8ddZBR952JG2uY0wYdSDImublWdmqQZd
bRLvLUD92jfZDkF7Of2qgj27EUyo5TEn9Xdq5scCrOUKq2sMMlTgHYNgtHwUfeeNufwPjC85AKS+
uzDqZ1bOGKTXByDUbuSHV2m3IcER2imrKUn5aWWnCGMyUSj2yr2sRBIRDHXhu34of1JzgF8GYE47
aC1HL7cdoNqCzMQIJd5hXNGlxKnj6ed6gnGELQwLu5CqsVLnSOISrEtENEsqvlgL8huxCFqpyEtR
/mDM04d7frFuBCVdS39bNiLS9Yii70FKpDhkEjT5k0+QvAXBmoHVJciheh2QoxeQ4p+253o1swfI
TLtp23fOD9p4aG4SRWOK7XhetHbtrUufJpb9LKvXYUVL7gGfOIw+7J0qRILeaIelY+SNFaXLGSG8
5TfOb5hcThnry/9A8u/Dae64koyD9rjhSy3yzpnnmauYFWkAbD0q6ofCeEGPlAdDMnFuwmfYjxGO
F3rdRTAHo/o6HfI7I7r+fdXl/rFW4fSbo2TxWAjfQm1wC0sFcFEp5yMU2LHSZr32r0rjyR9BSpdV
e/n2M0hoc+1sgFS4ykm5f6Wn61bvyO5MscPbU7XHOvsQNxDSedwCPyRBseKMgNwf1B8F0Ru3Uwcu
0tE0B49GWDkUfPDgX+O2iOJIo9qZVbgeDENfZ7CZ8ojKbd8svTlE0LTRIbmeVspyLDVtTrLPr0EU
YjrvlbxzuTpw9XpaFqa+XSCxdcdIpQ7VZEfueFYj6PrUmLuDm6OXPzsNvLnGlRVDBuLhCzv+yJ8x
ucubqpnzRbYaYzl1EOoJvM0HQnycMjkSG+IN6Z1ixIb/1269nnvVf1yHCZmjJrpuBsXBmMfi0SVV
ZhtCeWPa/Lh1EVYTC8ghQMGKsHgDaRm3n84XN0y9ZYj6G8qWPzl21qSLdUoX2v57TfCOHijS7fBY
Ju73QnG6pAF/aakz7uKADlsMcbMwS3cZwFv+nobvPYBduZt2ScZtjtNptyKp2HVW5wMeT4c6sIR2
KM5R+/r5/O/MT1htocevr5zvkt+yzVmEl9c7GKlScRrIovIhmba1h9x+8rGuf4zsUdeIH8B8q12q
yn5otHzhlBEIPGYUgWSJ8IbjvPsW6u8r/Azv0hhJ9l6wTORptFPIcDwqUPi7/9JDJk+aIrCDI1cw
8SVnk/EZ582SLMZZ+gM0fURckyLD559xOYzB59fa5L/URUqKPdt1QxIZZB4cNzBGMKLa7s3ReJCC
1zMQPoP90T/+fgTONIqwuvF10PXSZ1XUJGO8CzXZG3gebXjsJEv8lvPsf4ptC6w8HHaPnqiJiXBe
CzQ4g64x1B7z7ZylqtCPLLIAqmFP/lIhU2uNQ0JfU8K1V9fXG5ANHCPKU9bL7HdKK5RgcYxrnNit
DR7WAs0t/M0d6nJV/Af8feTDP7OV5sxN8hyWNGwJ8rOAry/4fO3aB0PX7pi0XJq20B+nkX25D/a/
G3jhV+6Kv3KiVv6whV/T+uO1Mdh4qK4Tp5dBMHJQMYvrakDkbV+7P5PtaJ7PrZj2UFjp/ob4gNi7
8Ex4AravlQ7bgwcG3cicngldALxIxQ9Q4blT35BACZf2ghBpjXni3dnFKBy9DkR1OS39KHw8WJBa
wymb33kPAjNKkdqajUy0dbfRPMpyxVtXk3wmfbtjq/jKeBbnOdLZN7QbOXpukzV44cMw6MArs+qM
4pcOEcXrWbRO98EdAsQ9aSWSUVA3uVGSfRYOSJZHO4gFYKDYRdCeTHCyz6bq0/7/Nzf/Z0URhl00
+vg4v5Hqb+RwNyixVllqs1lC2/4aClyO0CBWEs7jWAdBj4HKoIbo1B2mVC9P004sLzXt2Hb/o1Ye
X4DfC+7+4OPi1i6FOoZRIskZH1vldziB5qpa9OS8D7zF+DrHPZLpXOzB7biuhSwHOmZzNZvF4oyB
YBYQonczPQGUILNIDbQiHHoRHqzTIQ5NY4S7fKXPa6O+HjVNwkYI6zMd1tUevhq1Rml7+p2u0juO
KwIQWQ+AQRcAWsEIOe5Dis+rAMsrShua5KZJpoiWkTvbO2ndM0FRQ4XQsKQ4HWPilfB3/jr8tcwa
MjYP8DQ3p6L9h9T9n18rp3Aiyx9meo5XaAXe6jcYKn8A2CdR/fCbkvlua9pz8Qb6to+h5j0TnicF
NoeYxMIg2Q+c5e8AXrtMLtqNwhxmaQE17kV/0f9exSBdxtgQdrD0qt7QlsHCxW4SheXYV8RSZBy9
vN3axX/3/0XVCSasOOVtf/e1ybPhuQE1AIVgdencMsL+JlH5WDXHjoEwRYBjo9QnTqJat3M9cNyU
P8/wbFCekJGOxyzVl2Ca1seg5omVriQV2/4AiVOyUReBzQC2Ek7Kke9avN5xjPZjug3hDssqNZBi
ojPGbd1Xr3ax+7t02kqTbTv7o4aBmf/gsDAGWm1D4L6MvloM9B84gnuZwUUEdjLkFl3q7j1843kG
kPmCfesR5IMg29U+yVVfyJS6WxsQHs6tZbwyXXuGw0ZqaPFXBe1jDU60EJHjhR9+dYlQEVqu5ZYS
hyOEnnFUbx4dK+cxkiJKw4V+leQ9D94A+/AyF9msHBIZNR5F7d1kfYq5UZBIp0yBFm+msdTKiDwq
XILya5vWctiDA36qIziSWFbFMbZ1dcJm2zGWQKNLcSdojlsPdeGzNW/6y1ClZu6LFz/wnIVaBkPw
cWf+Sz+/Dqq+gNBpE8Fu1G8RedCbg8vopV8I7KgOzQ4N5VUYZDKDZLVS/Cw/koYtcM5sjNKuMg+v
uIiNehF5Pbry5t1xLgFDE9B1SdY0G3KqEaSX2njlogLnzcwj/AeFrGXKxjrTI3oqnqfh06mCCUto
zBUBxNQSqF6d3+LxIvHQGdQNQrwBZS8XyNAG3AB6sfEGjvrmwUVCbnoJoyPzFXMSxE18nKtnOeDp
QgaVIEs0SDAhkg84kaR5DPzQ3KMm2+7Qa/VltTrS2RABSaOvQim3RbORpWiHWhln1GaZhztsrP98
otJ0TUUNHlslf5sdPaiuWdFgE4VaGaOO0bAvY6KYXcQ3jPntj2pO7Df8Ssum/AWY+MgoxkNM3qa6
pfrPIT88sdQjFcbjW63QLhCkEZ0698PI0Dotig3Nijf0jpqIemXuj9c8n+ABXUVxYyDGkeCGGR3k
XqdcEfbwk8ca/+ivF57Q7+xybV6OX9Ryqy0fS3ZrHzt4K70+LbreO33ie+XnhLZH4mSkrAXbwxWj
cKDXDxYmUr2UMMPqmFr0jc9DSG5YaHB8tsuXwd+vXx6p9PL/+bBteIVbMh3xnsJyEN+fV814NcOf
FTZQ49DDYKTsjO9WKmM7RS1exWugq2DT6aw1dldf8a2NzjfpVQvStvrPStGdTrOTTo3jvMISjKLI
2k1qdw4zq11I8qriFavGZZBpullCAozMLJCGrMS9yZRlE9Yn6JNUoSx5gSjyPpTS3JMs5tP0Mwfy
gUno9LhqQ+ystTCy9n5eBa4/yqUjQ7cOF6rBcRv1+HJpiUulQgC5AtFIOxbBUVmENG8XJpJKEkQx
3yQZcaNLvNGFkt65cjzZJHU6o6OKQokr9aGLNzLW//HU0tlFtLKeMsS5x94sG1LhJk5cZ9QHqLMv
A1/alwGq78YieAuRhIXFoFBqD4fOsCeic4xKERUT7N9ByyfvNmuY40TqY2NLgf5+zKvbUt9Vxzy3
VyruSo43EcUhb8fat97Hi8AtM+D8Zu5gPcDLxZzexqQ8p/Qcff3COhBlqPZPjqUg6Xi2Mi/7Kz2u
Po92gHc0YaTii9nLzWwlrameHn955vgueYKe34yYoSM3Sa/Izpfk7K2228L/YzIsA/v6UgtD1EUv
/VUEId+tGEV9Wb0coJ94ko+az9sOfKvf0I49rP6/p4Y6nz8ucAZPr4QdADlXWQBetCTD5mcKl7lj
Sf4NKlIyKPYroeCJBpn4nIuoFrHOrInzhERnrUEMmC/BXsyCB14JQovr/PzlYmduuZuHk8VzjCRS
pwCVeuDqtzD5oHh4KHZlL39zLlQ7EPBHJS0GAkVqrmTYhBLk0gpQLkmvCE7vUcng9pgRtDCESe1G
FB513nGZ0yqj/QSxkeRNoSr8QuW/hkNwFgJa4sJA2lcGQ0VPdnCBnZ4JsRdduS9+JjQbj3MNahhj
6a4kV/WKi2DtlWfcom1vVobKMtCvPAa+6tPPv3mzDL86aiIK9uu/zNC1PfgidyQ5ZjejdBXvbX/f
4Xa6vKpOo1ikNdZE9LlsNjdJegMEyq/ypjxpCErTawvcB6liy08fYthsQ0ldNL+Z4lf+v/476zrZ
4LI0ZYQpSuTgyXaVoX6szDg0cWxcIEZTCZEGg3uTC4gGZ+YBeNx6dLWDZGUjUtDx83tUJxMCrJzD
e8dleIHhKncnDKHzQLRxox0ob3C+gu09jrx6Rp+kc1NxfbvxzEZ33uqtQ+MwJeHW+I1u7AGyi78o
wUpzTjNBXaBGq2halxhp4yz4P8oNDZSTDOVYas6SJqkzZzmvjoOG+zo4PY7mYw0gTl4/HzkeEwOV
rbDogGMIXgU33VqbHnnOoUufYhXkBjUUfkvggbFWwlk0LoMNo1jCgCxX8bmL/y4Ye/H8aCN1lJD6
Z5IHzIgdpOVIHEvSgLalvykdwTFqUrdmhALnVEdykjVWMO6RayeSP0Z/nM86lKY5fX8jbkOMNkpY
8oF5p+fI7LvXKfvBlmRd66+RM0INQRDYSmMUMhJm3eRW89Ok4IiPplKK2ugG4uvYQbEQNtibMtNU
uYBKMrOzVMHKXXgRJhixX1qHHqO7mV128cyD3WZrBHeFU1kgmrPtQqSGQCGUMukUDRGs1kBgptYw
lBQB7JFpcfPE1intPQq9LYx0aW3FcdUemhGNvk09PG9hs9X6IVNTmczMz/cfl1KubKhAC56EWuwO
Yw46qrgCW9VlduuZgCFl4ne4evwgSo/Sa/s4oZ/hTtaDMfu/YyYRUbS0qJ3Pz5TfjcH+4nOFuqVJ
aibaHaeQQP66c6rQvDs2cPLvpFf49MexdAqYx0pBttYK+zi50hAYhWGB+a8NAtKYAfAFXAIUF9aq
UEFcqcyHq0JEdY2kQlh2iGzSN8+ryc5BKB2NFl+rXqUdUeDQ/P9/wWzzDocEN32chhsie09TDfVa
AtkpiPiPI+2aCRFQ6CTB1q4HyYffgTq7mA8zuLARBr/fwcbbHXYdqF4GClHbxyUhW4aLfu5oOHp9
NkqKnTxjXbWrGA6MqphD4HncZcfqKABaVjMkhot4NrQH8yO+sUlHC+/drBHtbepgxfL/46/GLkgu
FKWQz1gbDbUOd50joyB58Gz+V7eneJjxL0/hR6MJhUHJw/JMXyAjS3zregYqjOWX3GTUiFCaqzU+
NdYMy529qnvnO7j+JsZopG5pJZOwkIfFk5ilhJEPDxi4jyeUulDuYlGElocl2ZZ/h8zP0GKWvzw+
wcliNXRTdIkdyeHB+eVw7cSKxA0BungsW7B6p5GsBEEfppDfkrHDfb7IfMeH4j0z20c/w/LkkG2S
JYlo3j6HurQlIITITt4zIjF/77wQdDGXkeyMX6B3gXhhsNrZHTQJaXVkSqwB9fxQ9vDG7lPlQBK4
zs/VTSWqCtLZGqlvsHhUxp70c37k3Qq19hM7gAO22Hrg3LpbOOejJzDjey8cEOmY42PTMmIxmICt
n8s/TzGhONoSFo+DDVAbbMDDK3V7A2nOPAA3vC2f65TcYUtEZyKRklzM3tjwoE/tLz1Htr2hmQE1
bKnUp4e+wuMztgAhjHq/XUPC5nUsJMhlCAvHXNQpZ1ksqQWib7yhTTv7QzaYm0Xw+UJhbDAveVr7
fyGhpVbkUbauDq1AifM6RYCezSewR8LwwwKVDcaWapEICcWk3eXonJoAs7FluApKNqFk+/4mheP0
qumuM6lyWf2uCxD0nMxC3qwU1DGAuO4q1hx6cZqKUTms/gD6dDI6A3XpTceJg3Pq0t4mP0Kf44d+
AIHleoT+KOh0Xez91fQxJWM9LXo1lG9hPNzsem9XPsTL1pddmvaDqqBQ/eIsv0QaClHeyAwAOYFP
lfihwKWJM/8ogerYkn9fVQGvCzm69/iJIRtPfechBKfA4w40MTAeAm1JKJZn5yCQTaEWZ/E7QmdR
Q50hJ68jZNN0L6tJtTUmN922MUmPSfe2ZWucA4acaAAcB5Dti2jxEjdiNxc4m/PN/TEiJbo5koj3
VDHm7Kl4Nz/RnbljkP9FGTZR4cCaAPl8GWP2PrMRjg7OIgmnpykMjgijUrI+0n1fTncdJrlsPXhZ
Gw7LPljnuEHs0x08TfkzHdHOoUG986TSyqaPR3NY0litZu/WGes838YE4y9ofP1ySZWubbd6XNAK
yAbfqRLJDY2lAqGjB+4/cFW0VAHspLUhDH4HU3FICC8L/hZgg9KFyGgsdkRZjF6PeSZi+3iBJHFR
4Q7/IttxgfV4deOIhD0DkSek9tmmTadZb1RQmBTaGgggzbeWW2QnhpVF+PeSezR8IEi5rwtQON5Z
sBnoJfKMZX7GF2N38HoAzcWpCh4HcqszvUOaJOvWk6ANeZi9AjFU2Acy2jqIZtrMO9T34gRN+Wqi
XC4VXfTXxaGh0CS8aSifhvFML2LnraV5MMmHZQq27q2VcFr0DSi6BYNf19aRiZAfoo1lL2iiyg+3
U5G6qIQRjZIGcqmxMKS2eDb+ciJk4uU9Z6a8oxCcm2yxevglBuNFA+EIZ4EHR5kvWhvkvmCTIgWZ
xXaiFcarDv0WY5yRgioN5i4doauiM4XW/0d5UPKT3TndRr9jODFXRgM2dDbTZxSgpsPMibStRKgC
hWBgIIWfy5BvGQBQRxm4I6OhzCEhyKimBRj6q6562lVDOw2V53H0P6VuqPdUTKlDZLJW3IryXf1b
8TWyfmL/1NLJYptZxEStre4iEIB2VOxYAmFkuhNl6KajNeGzBmG5mVYyWIL6Cqx2pYjkOQohuSLy
tZ+DnOAlhf+y8qmIyGPaHveY1Fs9QSUGxnn08FgvRKQWJDlTpKIWFKCLCpSpJbvrFVa6YU+5eKqL
U4VEX1pLdJK9dl+HBA6UFxonPHzTiY+ejWT5U5t6LrWNegwZzJzCwpBwxb9NZdPJ6XZaW1uJQFfo
TngEfwm2tWekG7PBMgrKjCqspm4VOqi5v7T0BCwJFhKtQBt5sqhNsl6Q9BA/J2vSGAosLv2BlSDF
2vjOqzDfM+5Nure30L74au98XlvrRrsLL9qzBUIlft4rp8kp2KEJfRLDTewy3tu33r/9nKWjw8iL
VBPhd5tjFBlTvTJoGzc09M7t7XNhug3GmFkH8DHRBC2G7CguQfBJzCFpxO6Bhbm2QpJ+xWRgQEaW
iV8/MXP8CoEX4lfygzX5IbJ1uboY9BXTKwFOqejIXHn5Dox5kFYg7edSnxVY0J1R5gZLgXLjWDaS
BuaW97vTQYS9Y6B1WzLGzVcTIOsKIJkzGBYk8KIBJNjVCcSgH81a4c1jEsAygyc3lqC0yF2p2nid
we5wuMjWJlaoIPZJK0TCDsd2UEsnrvMU4SqrMbphmw2ouiIFksKvnn4lUr4EvwOrcY5ZUnH84Akt
FqradwVETQhkHe1Mp5c2qp+nfdcn4sqEEGiCJGyTNSktyvlEkBHghLTXZ7qywSOcNc/58pxl7VPd
GUSQSCH4+xX914xjJoHJv87Ui5HcyY3FcqBnwS3ALXL4HbBjRZD2PcFL17154i52FCKl8NV9IR1P
S//tM4A2tgq1c1MhaqqURguxrk9Qtf32pXVhr04f7KG7dHFhaAfesIpxpdmneorwi+LNslQOz+UP
24F5tWS7SEq21R0DYhSShgsnYR+/fFpp9Q5mgEacc3vxXoucKQJ8NCWZP4Cd1ODQPZCk0tyUeec0
scYY3IqJ9Etx3REKGqNG9fuogsPtL4pLx7U3QP3CjyDk/80jmFKJ5QjRHaxAg5tTw8SmNwapnaiD
ssiskXKp1bt/L9DWPGyxz7v8q0cxy+IwbEOyuWghDvRHhb/GCKchkHiHIPvm9t3cjOjAkcylkc+E
Z6npyifnMM4icSdcy5fBvOXNFn/bTqPbsjGRRVwUV59GYqTa6d1J9qHT8jka9uPz02qSLWbUpxcO
GyQPNHcGnxMSkXNUF4zd379ulSiNKvrU1pBPEFjT13noezEmWb+A9xk8wdwcLOKo98aI9YR/Opfa
FCebmrGxcEpBZyI/0fHIQS5RhYRA9Eaz1qGunX4tSVqVLdSL3rHbyvwaDY+7ucAdu4FUkhpbv8om
K7CAXtOErSGWrXXtff/MQlcnz3fD+MHdDNm1wukk/k4zd1AsGVTVz/n5UuUnpX+xfmJDNulB3OL9
+dPfAjBgV49m3P9Jy7BVkJVyBuoHPa1/mBTDG85LmE0pNOpvDWqzNnYsmmbL2/EfTQIBi0qi3Ss1
TGeabJV6sOwX02DCbkJ8TZ7RjYaARpT2yoXBZ+y1ESh+Vz6Ya3TQhLiJTBMOVOSNkyyx4IXMW+Xj
vxZ0H61Q3J8s8Zvj9VlzEDm0FeGYMDX8JBzwQdAcnH51s+xc0rGSZY4JlhQfjUSL5siO7231l/dX
npHjfYNmp4umk/SLIUcuu5y3HHDpACQIRkYHCcNj4uRjyeQJs7soLAL2MW6AhEXMs/qN+btVTh5X
t4m16idzr6UPdOxDWBWSUO2H3Zs9eCLhoWYsLF4iEJ275qaMLgXFB6CAFGum206av4dPRzkOKimF
+yrLs7m6MolNOfm3eXgG502mt4hzb+9i0YZApzms7QjbFI21kcjScWYR8XGXPrbK7P3s1QCkmHHz
JLPXKOBzhmPUHqeRRdmM5axbFhjX1wbFGB2vSYHVP/IoZPbrZd1pAKZRD6bXAnhxv6Yxvg/gzaeG
r2RujtQIH6wSQEfaMjU4mp459MWiJprdQHTZlwy2nnIV6Tpxy2q/X6vgpRYcAUbn5yIKmMSFVtdi
q2pVyu7QWfhZHnr7LteUzDmug5G+4vn+R3FD1RLcoVYSl0l90BtGeR0LuA1D1nLKuK+xfG5hCJaT
U9Rl/Anqg8xkJ+FDE1pOI4RcxBN4nquSFosyWB94S4uZf9Q9eKExasGsIs+9CPKlA5EokfljakHy
btAXN9mYqRUE/oizztYtQqWowJY0BszGZK39lqVQoj88ageDtkGuRVZ/pZ8y+BpvG9NSIq718fS3
sQXtUhYk+INuSJT/HrmAv8WaNjOPBPsw2UwoHc+XNhSDpKRBt+rIHOL6KjErrV/VGyu0igMHTLsP
FmYJVc2tsJG/0wDAsN7w+TBjyjivKZ6i3sSsf67AvXI3s5D8CL2ksGbDSr1Hasnj5MrP018kKAdg
pdQxF4LbLhVvPYV+1GF/05u2XhL+C1lBaryVMDhMp4vfjDBqZEPNsCbpNUxCXjkElAg2yjCXT9ij
PJEQ+taLlXS/pMT7ZQ3c7gDcAbK1ITKmZGjyrv9S1hB+WA+VOUL8JC7Vuet4ePTZfjOzb/iGQVu1
W4b0M/G9mD8ZM8znNpWzonpdmN8iOfOmLX0KpQHfOg+hUBT7bxeKR+DtIfM/qE+iV4Ub/LDVDsYv
/TTd8XdIkAwGfl/Z9ouHt8HIj9XaiS0ph1ZZfcgc9y9lQCWBo76YbeCPXShY+v2lzkV7pmEOnDEc
dNtK9iL7uZvaz3hR/TeIv1S/Oq2Zdq8esDnrPxiVCz5MxBmZBPU2YwD7svVcBlmAPQ9CAZ1I4r1s
Lx1IPdxbHFnU88xY8SFrZjRlGaBrYxZIxb9OX2sfciAGwhm2NSiaxroywg2YFjtTagPWteE4LJeH
jpvCWg4PhRXZ5WQkhwL1INn9rIOe/2vbmo8v+mnRx5JuK0qRbqAVuznUnoFuS8LjMj9bv6vq6R0s
yA+pNiiopYV78sPRaraNRnX1xmkeiGlO74w6DcSt05hCVxKeCWhg2L4ZH/0y9Lm6flgjbjxAHBnj
eCfLiO0rR2Zgv8i+x2VQhrr0RpPMTeVT6QbiuZGowxdvsNtF9r0arUKUV0phAdcnbHaDLmIMB239
LbdG/oXxtEENjxQ65e5kp6wCFJNrG+Vh+Dm18CYN9kHCN3z3KjG1xdsVVrNmjP36938IsKvzKxKE
pUEGiZd0oWgI7n9tZ6ennP5IY6gufqeyXJVGeXfL+vcYp3J3rKSNvyJH0dtQTHcDacgExMkNJhQQ
PUByELgM387QavDl/93+18OWiJEKswMdcWymWuU4tBcQBxLoB19B7PXlrxeg2QN9U72ZzzM5JEBJ
ONlnDe2cTn2jMN1eXYO7rWLEt25pgAl7C79NQlyhK5ul3Gm1dhO2CL4FdUC5JYfC9YDFsWWOHLE3
pTTSaRA5sD2Ek+XUtVqYJ269iz+o2d2F+XnlJD8f/IQS8iyLv36TErRKB5WrLMpTFhekEA9OhN0x
loqhvfTDpJAzG3WWCyYQcM5QUol2jx8ZQYzHrKNtdwZv2R27zVdcwLR8uOG1me2tO4QVeEJ/3PkJ
30qKu/zQyFuKaWJRPOYLV3KfU3Arv60DaB53V7sAFyEckshjFmyTE1WOhDnRvouZAl/MOmFXFnJ8
UtVGnHGU4Y9FjcqdPWfAGYCc4mjOr9AQM6XcumLfBPy5bi17UAKPWMqTWA8B4VHrmnx5OO5/7Vkb
RCsyTEmfT84LMYZ5qSOpnYxHuIb35wQxoPsofNMXGPjayL5TfamlZyTVLAQhS6zSja79iLw8teFr
zbQPDsdVTweuVuqE7AodyD+pskRdErQjL3KCyCr1E0kVKvwxJfgF5glYCn8bVI5h/3V0QzvLKtc0
IgoGRBGx6sXyvit+R59VWGDc8NQotdVrNgPrOwwuC8/ebYn5/VZV6P7+DwJjEAPh0a4cgPZ/xQP3
DTTVm1YFUBAF35OjxGlZth+dJe9UtdXx4phf8add0ND/4X3I/Z4Hk1UoIc/4aaibt3HwaqzupFDx
F22SjnBkiT92UqvUnwb5S+FFHbrQTGMsuukuCDvMTj5ypWYC6p0D8vOQHBG1vxwscE4qRSVxoY+I
tyVLXzZgN5tAIgkQXmUQh97WO1kWRM+6SoBewp5Hsu5JoJyCukrPEA2yclncFW8/myi0xWNH7laP
nNkbqvUbYDA6k4a8JSrSYGS/KVn7mL9oWFRS/MT5j/CQNXTRk16e5/PHgCEvVwhqthb2est7UVJ5
uwvGaX+wMsESgxu1IiulYGAigNRfIVo2W1Xou8IiNTP7QUphiNljc/THqtRclskoizoyRil4Nqv8
7UIivk/6h8lCONfp71X7pr2asNCy6Yjlt63+NgAAtZgIubruBJCtHsfe2lZcOf5XTAJXHvy5lifJ
SPRYVSYNua476zYJKm+aL9ktB9Ec6clJNGx+3QlmUhKC7pghZF7aGUsfcg51BgCkZuerL0ByGkuE
qqj37NtHnY0x49Xp3xT/tvp0geu97TqHIFlXH6lGDEzJTMoYjBgaaZH4F8ZBWLa+zI9nabPjo9WB
dK1/aTtBNNy5Ig/4go86LFS7YPrY9y8PkzwYcCrFXi7dLijNnb3A9H8I6O4aWqvaoAsxSMj6Mcvg
PgjHpLwhmuC58i++dytIWAIq+lOx6qGkQTuPaSzgydubnW+Vufat5TtS6iwohzZEIsVy1uH7FTsa
MmKnyKGFVY+ZJosifWmj/59iKaYe7LZY/khr3U4TbWYsckQw58gbSRo397nipxm8dHUu7hNC+09H
/Qze12rCLZkv7kx+9pdHWUJ6QIFk2MsrEz3jzoazMOn+A71yOOy+oy1705VX05gwdpIlin67Xiz6
NKcXQugAmNYf2QIWymXgG0DC4Y/xiA98JGjm21mwsQoXmZ3520y85SghJOe6ocXh3c46j6Y1gGLi
CCPPWXyJKmXvwPsJE0tiXEJYIouq8poC9LnXBedSA3eOeGCvyVqlcCt9j74SuYQ2F3r0E7x78jAx
DRRTyp6/x5DbLpCeELyIoJ9z2yZQ+6BZPzCjpOm8FVW9j2+C1IX71aQTM5JD4tT3a3uAaZ0q6VYJ
ceHrOgOMR8fwCKQyDlZQ3UzmzAlZp7VKx3s5mJKPFqP+yY9wSdAjmUHjzNxpMQ6cF01JynsisBCc
wGs7jTPzXALHmGYiUQ2aH9jIhtLFrVvS2VcksupfbyWkle9LXEFxVLAOY3nBw9jAWoqWuMk1Y9LF
KFU9APdcVet3GncSh/WGz8cK7bpecpUuIhZ0b4NgnwfSVh+AwbidzzRpEz398RcJdBHQ52olPLJh
wH4vTq71mlthqjUbpQhEBptJf4j6i1BS0sC12v+awIk5sg9ZwS4jErg1wrh9IVtt9n5kN1Cu9io1
rkiAcO7sbJivm7nfdgLBOgE3mEmrUUGbfXdbCRKOYhwD+IQ/nLbt48E4bKR6m3MjRmO7xaI2x8OA
EqiqMmL6PhMcYf7ujtxZT9yI3/OghN3S4duFznZsbQSVzwzEKmuHl4cLbaMgm7pjtYPyQ5Zk2LYD
PcMt6+0abTalYOtV6eDcf4Xh4SM4/O2/GUGcJtaDyhQ36d8HjbbzQmQK/u92YPT4SH5518dZVREE
rnN5/E0c+csEanNHfpKOLyeLB/ek2Zgut8UltWBtL8Phu0/S9+6lPrI/PmzobHa6kp4GQV66MNiS
ihL0C6a0GlzFSDSKIRxcZ2rUcmN50ojjQpjpDIHY0kGdc7Lvhfj9gm8XKcZKK8f1d5SB9E0QeQLc
KX7V5QzDHCuuad2ThfSQIXrEukL8NDCKm2bKD3z4I4GhpYMWLL//XKYgFLzOfGHfQQLspqlhYVfE
GQjHN6NzrxI0Ho3RdzRRhniN+pBYThnxQabtZWMOEF9lLYS+6P3eCxjpozt/QAppU+FGccnxeMr0
0qDCPpZ2Ie2GPo47AGX+kggVqMCpn9jOG6MHZL9B4ztstkoujlkmkwuawMiWwQQOmjDM34O2T9Z+
3gv6wWBYEYy4ByKea1WtlWToUOZexX0vJv/RufFBeI7FtbCaY2SWHqfGUItiQNhSvGAyseemvnNq
ZSTL9qAIkgBgdva65iXrgFE9KSa8D6Da6r4cimclABHo9uNFCAvljqw1CdIadb3JtR/cqdQA5n7X
zsaRbdDQDcz6PymmwEdtswW3EHiJWZaIjijUgfITzPuFHkwS5MG0v+8w7vyP55UvWpFeIrk6cZtV
IFOSTBO3JAggPuolit6HacLDqUYA8lDh35cunrcNuFOjGhYvfl6IYcJ4f+7iykiTO5/vQL7yZrku
nqwFE8PFZHZSLDL2FrIheCTJC9UdCIlUXP1yjgbGI8ixsgJtSShvoXHQE6mc6LivsbJPLbzTj1qQ
yWVB2BqqC6/egzE0mkjikUhpYIUJnvmO5+M20Ew46lifHPfGT0NT9LUx478h/K9fIb64U+505vTg
cjpkqBGStRCheWZxxlssNHQG1rqaCJxJvBJ+8RXTx28B76BFXthZc9MFchCs1I7BB9mbDoCtaqK5
ReWrhoQ1iPADmWWW6gTTqZcYnwqV5gm7VKPmT+EThiHW8WZxpwRLHr39mreUw1vccBdIygl90hHf
eaYUFAOY6RgPoYQU5VIh9zqk0NBr0zbXKbPpnTZYdRDZ033WvmeUOjpKQOHB9hlDFXYW8etN1O5F
hFiXtruNybUwQ9csqDQq+VXQ28SHNEwtIk9g61vHE55RLiPWpQI7ldRLQ8nn7GEozUrXDiNH9O08
Ub3dGdS4WXarkRK7kzr8bF9xGMFfidMNOOab0QVKI3wcGDQIvbbLdA8oHY75vJT925DgKtH8cMei
XtKK7j9yLYupa4DZE6tB7caMCkiQTLeKQYHyyxJ6i4vir/gn0unvaTagDCHRCngOHTypvHq5lyK4
U/Zk7S82+HvGg49/lcWoc/pF68wOwgGjDE/zHta6RfhwHjVv+px/ojJZuyxeEJJB5lPeENulI8Vv
4EpKeDLTIYnqAMqlE9UQFSukW0P/zWxONZVkcF1Vlcn8DzLUlP0oM0RJaHskrvYUn2nkvOe9KQP5
yoVW34niIKit5h7fL01dZVEBNQegih3jino6IEQOzpH+pLePSdWJlMdBYzXBksSyXIu8EVmQny+5
NevP/hKogSQDcJjwjn1CSr4umWSG6nJ7BuaAyqWbIFeImnHlByp4ws8m1+D3xeqn2CzGUUzk8bn5
1JycJqYxL/xs9rOcUIyen6qxsZ1io4zp+1FkgIm9w2ACQzHF67XOJ2wItqMS8QnisOgjEVqe0uT8
+eWbkTo+RgqJeQtY+17mThbkDeDAMfye2x5p4Bc7jK2Std+ZEPRDcv/f1rAbhMpSnyab8yBx8Eyf
jR/PhDBAOqClp2EApxIeH6qfzF51E2Lie2Wzu+Pw9EW9WnYcxS72ZI4KxoW7BypagyuV1rBfZmAq
SKgvwFwcwmlIhn8+3O3DDfGF0IIzI03ve0Y71GPzZckk9XWZ2QGeTxeuF1U6c4zt8IyUA1i5MQ/f
gDPevrhOPo4EokSLdXAXSvXyiTNpL8n6PJ8hq1WLBr+ll2o3yWjOVUzfGl/Ge9H4guNivbEpvuup
D9NeICW8OqEBv3Cuo/kpOB7JmxB4vl/8Lm3JngXKaSbYNsJtegCELDR3WQsiVOWmwKOSbq4vbknE
X14BOYOL0s+4uiqY8bgschd1PmXfEfCqJGjFlx6qc38XYH92W8thnbePnwcSEQLYwIJB2MunFsLT
Czmu0d0k1s82eISjihir0R3H5MXI42RpwFVkzNojdiANQ38YOS1zQM96XWhTwSTxIheSS2nCmg37
KIN4dXRbji6cnhi2+Tu+3xp49adem0hXDwcSGxamCzIxLkZzHd5ZODGs43HoCgglzXvqk/ye5ikR
T3EkQ9qphIS/Ng6Xa6PVKfmBQc/tDXQO4TWphBeA/ucgUG3kbKmLc196SFqFtI0EPfr1BsxTWTp0
q23UlPqxfXS4TkmzC0ZWTC/kdjmm12FaMzD4XYcg0cBf6DPxv1jPWIV8ljnnAiVm4iu/HS0MblUL
CUlKgrFPlHIgUdYjF8mAH03j3z6yzPbSt1saIRA9YNmWUypR6kozbB7qTKcBYcOqmTfkHA5iXZub
9y7ceHig/P432183C1qN0WK2T5QA94d6SIWL/rce2+E1Vg/XrGhD+Qfvi2lGXD2f3wZbKGvvJ1VU
IGzzFYkiYrA+O1/822ZjOmkI+dB7t08dNrUx7xj1Vu9jo7eJOcLlfOGTMrfVad8mK1hmhvIQBDhE
cZTPkUJ4Rno8EbEh8/0eiz4eK+AkiNV5/pOyPH2tTE8KsFCskxaJdKXDxFMS5g3LjV1J+SgeiXcz
phHcwn1tjlXwvepoWnBhSwCqUZxJqYc05upiuwlkZRcy3+kEfB91WanTe7wigIOKDDfP9McodcNp
7+2mQVE0+SM1RT1cn42SRgC/TNxfqQwwxvSScSWUhqLFFCqPcfovS6ZGmaShx9rB5eBkFLhOhSSa
sWtSGGu2Ot6bYsh0LsbpRrH4ieotMjNBXQLyqkKlx1DQjNBtVLrp0K4pRxr0AYSCa/5YIJF/ZDaN
jlrrWS8vSMXGL+Uo5J79MmH7Pf9b0JJ8lmzbTHk+OEpWSpcA0cv1I/vcxa3LGCIL6Zs3vdtLjXJh
M9RZAjoL0oOEaLYOmcn4P3B1FxO7u1atmmofcGEX5KUb38eYIRL28QTlgvX9gNDSwNP9DsuUvBfb
hkWc1IJt8kENcZZBR0tjvzgpD3+luywU9uqFZrwwQskHIrgS73tD6i9JZBnxIz0oOHUKkNxmQnry
hquURwcvxRkvI+H1uCcll8cpoFwRETO5Tm53b11b9W/nav6ps6RO3t3QOddFyweblz4O4Z33ALyR
xdDv46jBBSYXPyhAhTTrXL6NEBXOYcRTW4hxtNT7G3vvBaYeQ35XzO7h3y9j2ynbFrs8KlQyiIJL
2L4L7cUnU6b/XqCZQYPV4imrDzY7JHglelcAYVnFc9jbaDUEaOC0bML5M+ncsX4lul3oSA27TMZD
AWZ0V5loXExiiPSBLxt1CzGwjjnGN4BRvCT86IAsY2J6QHAtja9TPWeu6zmJAsbcEaoxDfCuL6nW
7kVE+f7xeIG7dYGcCIZ/yq5UuIT/iupSsme1A20WoqxH/5hO/Z2ULgaxMc4u8cAO9ufJ3J0Do6Wd
anTqKCXkruL7PWe034yUade4couLsmm+INtscuzva3FmNdmrWmcmsP8SphLlFSNNu/K8spVFdhHV
3dtGVh4zVh3ECKDYvR3MH5A7kwRfi3Zx/aDQj03jSRUJdjHF98gvDRZR0Bl0kjN7qVawwnZp/AGL
ulSp6f5ooN99c3t8772khk+/yiJYP+K9ahcib44NkstHJYIDPSstIO/3FDklHgifiYiDn+C4BzS7
kMgmfI/Q/SnW6qBhq3gT6bHXEwNNhB+Oe3ryBd7u/cWSKFukuilumFVruWBGrjkwnPv3nzePYFRZ
ODytM4pcdvybNEIYbFKFC5ZyaY1gyr6RECnbnEh9t2XQwPYBlfDNX/yuqA9WwtIq4oCZP82RrkzW
O1vn9DBUs1rwCbKAw9qfGDebQD5oHC2OGv5BOBg4lkYNjzjGsbSfKhD9q6tKKkAHDqMYRyvPav75
jR3VvHgIwmBM1cMXnnvQkMGBKJx28Lb66ncmi2D6RRXawIq5TPcsA5BNmbKJDxxHXR9m3yjKgEIG
of9QATfTWyFcicpCALSqAe6Q5pBqQuxWq8/v1xKEGPmaDgXYBczGdefUnR0VVGU/jNbPCgfCF/TC
yj9PWOoJYwCJ6aqYc7S3N5F+TtAcBYn0zNSFU/yoknSWUtB7zYrCbFRvc4v84e4EpIQJbDtota1u
m3Ll2SfFBAlkXtpCA12dFn0Wev/lRFEaO1hnk0YlyasmVa+lvt11m7CtywlVFBgpNXC+aYL5Rwgx
lnTlbb0QB8DmNi1DkM9ELV8BwrxvUn/CwXIjGkcuf0VVnDIhrZOdTz7E9wr05r8VZVlAWjVifGxj
qF4WOvdUew5zugFHvsCVC5uV+gkqh0+laeM19YTfmKbxwiq9DaKAGJI5Jr51rLtrK60ztXcJK5wt
zwMUMNYnJ8UsOnkxFISLxOFwEjbRdLp/ZTCSuGGqZUD1qmzd4JJqqEL0gEcy1E3ID2S2iPcrReJQ
lYHnyiVKmkpaEphJWiwsGyA39BcUzOaYPzzWHprgpmTxsDoX+DofkLW408G5Xj6KtbwDutbUOwjp
jI87QZBXCetMYGtixXHf88by6luXQ9/OcZ+8vUf8q0LG8JZf+pvF2ME5Ft2viUzT9e9R1oYVqHmO
v/W82Z33zc1w8249+4CMpnbimQ0D7+tmNJnQGppc0+6bB+au+2/Y7rD4ODPEX2aGCnym8H0UkfGn
6hmDwqtGDM2Qn7nAnzv5Va3jXjx1FDDx5d4uQt/jXGEbsdMB1rdJKZPSQpxQaIywaUnlVlqtV0M+
Fm+LiDVCxtIDC+T7P9JdiEPiRAuYDQLUKNqGwla3LIcc6FezhvkI/1VdzrJ/6IuW5mWAfse9H/YC
Zzcnf23QnXvWaW9uHhXP2rQSp2BR1LbINNf6uwnTerLrps39KLzAteRkGBWX9daiumtf2/ps7mhC
3IIg6Tdzgz/eVrN3kTKAl7uUp/UHC7TEL+Pd9RlzxhvniMCNi5daK7mSE9T3/IsyFp/aqsJcHtrn
aHdAy9d/JqO40s59N+UDnyAA9Ys9u8UkS7tz0l5sIhM6l2trCy51b72RrjmmOY4zuHrbyEc66BI+
RiwqP7J/HjXhDjVu7JTTco0IKad7HM40tbKMqVXux6r6kv8DqlleJvViD/keoX0MrO+0+JDhpOUW
RZTAbzh0DWV64i6imrGuelPdtwr2LoBQ3IIHwu01SxVknzKjX9xSiztrlyLYc7dyXvIU2WgmmSaQ
s5e7Ic1pwxOu69FXrnFMtbgTMhUQYfmnIEzx8ANzGVqhT2Bkfo4dY/SmA55Tyn7OsAviId9dKWg+
aFeofDfWNOwT3tbfhoOEqI8+oQ91Vem6afX1euSZsJJ69SvJzRlDQSJYL1DIMt8OdbN2oV45ench
GXxyJcuTrRzQhu/AVMitMTNLf2tzFPeD91TMyP7f43Xd/JopS3FoVsMSgfTypJFeOVqKec/vbdGB
maGvaRxm8rBrW51h7hp/e7Ds1vYBwls+04SpwVen/YhFMqoLc/BudqhfnCCOiqTD8niodx3JLg4Y
cVt0KarAAh3GRLGHzOZQgH0IltEJLLJ9Fe5vL0ACSP6DeeMN4VkrUi3LXGAnJOoBLJgtpqoH9m7c
7mjaqXNDpPRLLWElIe0Rf6XL40BfqGpUoX0rug2koCUj4t+ph4Ec/656Tf80BX+BOA9sUXxWJV6A
r3q+pnRS2Q4EvAZ213ZEv/uO+NPkluq6BeYA2XzHIXL//OzLcjxPUoyc0hCTUBSbT/eU/JvZx7U8
qYX7NnAX5Lv+AMdKp8Tc1XtCSdprMJbtLNgmW9rxqIeBCktlQagzIuWGS4ETdxUAsuEJnMZTkC6N
BNNPdyYg56Wq95kgHkrQui3Hf+wmPTxVJOXKDwncbGkskV1g0sm8QiUUiZtx5aM7z7JjCok6h8sD
leWw19WPFd12vcdpginioTIm6+d6HM6RXIPiNxwQEyvrTnOLaTXgWm5JCHbxs2QMaIEKNQdVE4UK
JaHv6zGmiYf4a/HpCyYwRihPTdkbJuUzaeGOBU8elCT8lDdeonS/xuMLKL+8epVl1VJldS+nKCr4
Kt2l9Tnc8eOmMXNKYJBYjUGQkfeb15pFL9vXlAt3hsDDuth1ud4eVKqSwENdh6KGZ9KRCJfO/pS9
0b2T0dFkzGQDCncXIyaVu1Pw9KtAgxAE7sSUa6UvIGxSH2bA7xQRFLdcHGEBRUy8KN9gXdkEBAl9
FDzedyeVtuY2pk1yespldflmVZwnR9RsF+ds2O25lu0uwhY8+Koi967Y5ciSWYfr1Gd9VbqDEMgt
GXvVHiKCmWIJzpFk5tvdKnMVS89wlB4rNUnretxU65Op4MEvpbbZcxeGi+4k5ZKJWfXt6ofV4iBz
DzS9MJPfzG+cRGva59P/AkTnZ/cRNwuIjh8X9gN1UmizQXA3k9CbsUWj6S0lJ+eEcDkyoUhrO8zD
t4m2M09P2jmATW+rAnKz55cgEAgfcDSANlignNc7adjn/nuhcUlwcgZ4iXD0tI+7W2swCXab3qLw
9zavO/T1v4gLKB5V34W+vAIwlQtqEVbLP27163KQB6xcJQkFyNLw5Jc9ZtmCohoHU7aNIjzFCQg2
z+/ZdE4hRkdpUeLK95em9OLPqcBHwlql9M3AcryQmKwtEl33VSCmQyAlSbxppB+KUSbRJK7hNc9M
Cqtqwp7s1V9ihPCQL06cC39wzYvF+iSBPx3aJKDZxSuQwRlZo1KSF5oNAQHQfmZsXlZwM7KYag8I
Lw/VVdrYckFl4pyfMa+tqBOpbQnjcXqXbtCjFwN6/huV2EPeZKDrBesq5PQqbCq2ekxSt1byaVHO
0VfWMPkPj1kvbWQnikfv1i+znhqdEMhOtpeuHYRcnLdDwvktELq1ohnk05DwKQ+HwWGVFWp4FWum
axTv5IVmQ/L1CcNMrGY9L+xWgDkR1bFd1b+UUESPsBH7j7EdmNMWlgPnCQaVUivpSPwkwR67yuPo
kj2taRu2JIwxmSp4JxSvfrbFSj/6zCrrHHj5h3rQwMmQwEjBhCe/rJ/lN0wgPnvEOeZ3RlOznMXW
NiJUHcpt1tJrWplLYtG/94vt16IdKRr+FCpPlbeaUg05HQCqP+z/YzZ1ztTy/HT9fGwz8hVXcH/k
r4b0vlxK+LVSIXwYtxuNEt94t1h5DVHhzd4v+iVwVrr70IAB9zRszodcvlPcsq9eA1oOFsz4OHE2
4XXrxHuJqAA2gYckLyslcyRKktFlVXNAASQj2zn+z+3m4wdtth6SGQwkC2xOvGUXhPCyj5SRuCdK
tQIl6KpWMt137AJWEKCE5//5QWx71BtPfoTBcDMS0T2nXVQ+ytZ6yvbmcxUPp+p1gAbx5Phh+uO1
p0m+tn69YKPbhuW4//42Picdtdb7e8oiOC2YSklbijSvxt0vZTBN+RwOo9s33qDweYGZMIYc8Kg0
QR+ho4eoPON4MhhYYYScuLUOfItznCK2MB6h9mkjiZZgX6u5TpJYAfSSsSV3lzcAkSH0y2VXFOu+
hsC5uu2mmIlALsREqOAEuF2b3iuFBmYjyBWEBLOmvS2JBAIDu5QatNpQtcZWFj2MHnkUmEE2zf93
/ZEVGu6fJkbHN3RmBUa+eO7Pgg6iQrR6zy75R866tWM8sFAmbONoraLE5yVC+DxcTtcjVrkuSK4+
+gdjG74fl9r0tTQJhrG1jH1BQ7XxetZjQbq6orbZUxP20s57bFtf+ZLfJLG65sAJFbU9c49gukmL
cwrUnPjOFH/OP/55AoVo7L+Qvp3swrGEA2yW+64cWh1a4tGc59qhTa4xsuR7rpyc700L415zaaWY
fZkZPEniIHtZkQE3g89TKS6CF+g7+xru+a5QCHWPmPIeAyAOMbdAG95fP9MRBvAiv1p5Dsy9oyG2
9K99F8ZH+GaaSMuOvEMnFr8PaKj1PwDU+NkkUtSAPgZKqGM8lGhSjNQwOUwIRFwFzBSaAlOZts5v
pb630fl+PTn7zAvqM+OCCCqep7ZTpEsOiHjW/IZ0q+M7OS5hnMC0j8lXIMYAw+IS7kKrCGy9nInp
OYwKQ3h46yJ0NKEAVfBZx+ztfmRCCR+pqyxjPxrfYPRodp1t+nMnw4iR6q57weKxbvCJEW//nYk+
1+GyA5FSd6aap6NKecIKBUTIVkYaZZRpES6lomaGGYqHTqoYxlgtY5bPKzEMO5ObsS4NtntxD9Ws
6K6Ylua8uya/3A9EKbOFnTcRf9xh5PVZl6RPxtFXNDDScq/n6VzLzV8fK39b3YWvih1mtQvSwrWZ
0JGOftwmQkiGX9oMBcGhPo3GubGUdlp5/gjvNuTK1MvzpnXJbf4jTK1jRdWPHGi6oiC5dB7nelhx
aHa+mRy+rtQu0Fv8QP6Agh00oR9jMRrYJv4k2po1nLpGTT6dCVYO+tg28L9+3MyEUUhD/iUiIHWt
fe6ONrbCSPuOE3AkOQDee9vsdT0/F9fdIhgD9HjrhUGwz4CQrY5XuOCIQweWATYCdT4R5Iw5jBzA
0RMG7zCT79j/EkoYd10FGfZPc3xGjPnRlUeJOeczL1AhGWgyiBHWaeXJki8JPq2jvZDQY3TzujgC
q9q6vsUc1TF9K09M8bz7LgVo1r69Mos37MJscgIbWBQvhuuOd1PpcbGHE0ddawtWQeYz5uU4KE04
Daz4UZ9budU59HNNrhJTU00kW8T3xZZS4GZG8UUise9XW8L4r0KXpgqtb6yRM1sk7dADpboxUU1j
0FBx9qnQbQO3U5j11cy34vVzchYYcrbS1tDLUpA/cSUGXtvaFyxJ9za3P/WcbRu5qTx6kPJ1VZXr
bzznomtzc1exrNfyg+AnFatWnAyLNpYr50fnRSjNHcDtwqbsmm7SbEILpJ+s3NgaO1R9Q3aGPFbY
TsdNvH0WU+pBlLKdTDg0YDjE+dRHUmdoGq1BtqoyGDkhkRZmP0LNac6dBiqeMWEz4Wf/hhrnaL/M
X/LFhoFuN+F9rM36QCpq6Nd5JI61JlRlxENl8t4t8jdiwsSdo1v5lEK7zW/zjd+kUjx+4NJIMxkK
rWyaUBRTsWdVe6XWkt6WyHQyOL+VXTb2aR+Fui4WIG9QXGacGNZ4J/JLpr58JV5/P4OZplE0/gh+
VBdv6ULTN0DWjzlNKs7ndfGhsLX3q8qkjpE20ZpIC2Vli9RS/asu9Ta0riZyA8FplvlPx/YNZgAS
uanGfqO2nIYGR+4gDFDyDPoG4rd/PmtBdM+a+cj2KBdSdy9JU62/wZNry9RGitj3YCl0zUvuCP8i
B7ehmTu0NGS/ADFsRkeCWkhUMe42Rn2YZf67aGwWI46W4x7iXQ3mrtKX7DfiLprGBlG6Lv/Ba5pm
M9LHGehVTy9BgDXi8VbQqJQDysm4YBvNsI3yvgAucGEI7xNVNtrq+zOULcylRez9gCCw2JDApUWl
Ycg5MR3myDPFV2qB0kluGIqpnn1nLRp5jP3U93LeB22zqHgZTwDS0iI3kbvB10ER1Ttb+i7nGzY9
sWc/r4S88k9m+PcE/ga8wJglhzBVuPOPrOyO1W4rE4K5xOmrHnoKnr8CmXd5N/cMqc0nE18tICec
uLIFSfN/bMMQGDDo6VCa3Bba87bAHmnBUpU5Yx71aXq/1OECWt5krORqiTKxoWX6GdsP7X14bfHh
XHnPhPZEGYwF1IAQXtlFPNpfwzoAS+MeD7XFx9RnEi3AqKHIRykYnoHh05SP152D4G4Zx1EISGyq
R4UR32C2JXU9NTULLjqe42q9ttjSvvpBK5OLXeRrS7mtP2gj2oNPUdMwPAltrS8tHIYP7PQap3E7
vsd6jpfQfGtaJC3DMhjhIMR6hADr4TJnNmDkfmYxFi8KyTSbQnm0zgKYaC4UFitmS2k+7jXzFu/l
f+MQLhrdWSpXsBUPn6z1VGxiFZ4wj4smBFZT2J0NW9NbuFSZIMXNubn+mY+GfNQHHH44TFHeNdre
/wi4mYuKdaXpyu/62ldGBuntj9xzqA72KgDHgzHzm1eRUQx8dL/PKz9BrIV4+O1gyZfqz1Rps22L
tdQ+4auKo9f2DzDMOad2XcdNRsMmjQieGzWTGzK9NkxE4L9mRC63K0jnqiXZ5HZ9wJcDVJr9uFeL
xqb2nMfqPJmtWOQ9nFjhjdTWwszA81gL6hPkSkbfmIGfljogm1rW+HhA7oCJAt+XG6D37hQtep1b
hgG9T96Jqs/eUQS7RGWpOOt0+x5u+Ff3FWWt+io8W5B3DE0+flhuyMeGLGX8iWGXgACLhUynNk68
rQPYFSw0GLfhFY9SZT2JCwWlHiX7VYqtHkJtGZeOxuw6Clauqt+I3Wz1J/ZNWiNeiZ5uB0dwc52t
i1/vxR5j7twyOZLoAdNas4lZ4MfrXkdrN4/aggGg/stiKAkr6FTFUCXXpsLkKZthCGIn1DQ0j2JT
jKiaiVweZRRHnjb8ZKInQeBbAH4ltltannxQt/1CKwvzjuWriJJGXES2hlKlZZSmswkuVJoPpJXB
+RBATNK6V3V344IM7RyyZbu6u56Bdc+ix37EOAqGZtXj5CH15bdSfCl+3X0aYz67lawPXsD4RzAo
Sm4wGxHNaM6vKS0h8bfDqUvHhIZ3e5snwA1o07mpTDTSL7ulbM53fbz9XSRijJSYhjXDwLJeA5nJ
tPaJ2ZV+9oEGK0ha+4XUCWBknl8oAka2e5x9RnH/dPuwYq0lMiHT65aC1nHa6JlBVWd3EAhn0Md9
5ya6mHoXooGL5ZHgGEC9tEAob0aG2mknjwqSza2ljBGIuQn7eGkTpG6SxuLx4eTZnN+SsDXP9r7N
2OISm8pTORSRtM2LMr7X9mHIur34nzzkfCkbqjNud171Ze35A/0SypUrYkFSyFoT0q/LfzDVI0Uu
Jt6+BBAcmBxn0Cx9BFHQW659iehIdb+WKp4KUizahjZAywW/a++z/KgNLoqYQbyUALwMrOqz7J23
qv5hxtoAfMK5OG3JgV8FF6qgjm+xdqX0hnVtap9kWGEeYTge+JKfKHjHxUU9HohfFgjeW38H2zUt
Iw+3Yrnzz1Ye+mlb1QvL7jmGRfyS+IIbX76lZyl4P10sppuI/ml5hNwO77BDXFti0uksKq2SP9zT
qvaaxwEWJQkI/zcZSlN9+rfyG9qWYw6tsvZZI3X9//jncSUy0F+oZaI0Y0IIyyCbLJkgCkH1KipU
0hlIg3f9qWSUUB2YF5JgOUJ2ZSebTr3ANFUBFWthZjwKU9iQbMMNtP5J6N2iYjhPPHcJcqpkSqyk
7sZC9CgY0Hgz8NTfcpB8Cg7inWTY4pUYaYWsV307guc+cCUPi31zicMAek9vlD/jGvWkIjtC7w99
JvKdQ2yg0mfdBR3Cq22h6qBWuLiujzRR53AeiQ5CE7v78fAt8J22+gsclVqEFxvcQQTaVvPDwcOJ
rqPJdUsbcGJ+SoR0iilrEF4hv1eNESPQPbDWnmvD/Q5jzGPQksrs3TIj8/Y/qDXonYgdbBAzTwml
+x8iV8h0u56pfRuPwaJAs0koGiniY7ZI2J6Q0FoPk7v6AEfrd3EiOI0iM6VPXLdsypzbqJpXvWwk
8y1dlNZ7EtwfuVdZ/YFOotK04lW/5OIDToTm7+pFJ6diBtIFyTEKH1S/YCKlZFh+BfvlZGQPNB3S
t60HMOx+u6XbqNEVb+QbD6PyEWeA1/C2l+l5jwMcMS4h9EtY08gXbDT0QqOxEOrqpeRK3kGFCd9D
RYWpNE4XYCOAYqg4MIijXK7NdsDhrHyow+gLFUdZnMIvdZRV3Hyi7X100NrBnHywRQMJ14Uj8ABK
ia+Dz17itNUnmOutY8oF/MrUiW/FOXH9CzL62HK206K9wg7FlprLsjEL14XwDLyFP7tBQjaS82Uu
kqrtOhk6DthweC94oH5f1/GUs46l6ThZtVvkHgjjEm6H3pjqaxTY9d+9MuHpuLydcpULS0iZY19z
/F++eUGfeyhJegLViINlM+jmXCwKMH+hmntB/jDkAfu59j9jhWK22GGJBbNuesZwoHP33fHksxKi
rOi1v+cgk5xuAs5G39CRiS8zaIKbeV0HVjH0KkPt+oJr6x7YhxyWoXFkVA1v114vykyAnhJWLLbU
pGBrGx7OV62O/CYPfaqqgcylHWOTSLvEltu+NGbo6Iue0zSW1bVAuQingQK9miHOFNPMoTfYIy+J
h+dV52k2JKcuw3/58TOrPa3O3KpAc3O6woItSI5iQR6sPW7Uclc4bME+XNzROiT7rbq6RAZ7uw+K
tjBUT26BTdOqFWv0JcuN4f2IFKMwKbud0ThSf9YTNRO6eNQtU8Hk9zXxILxvOOU7UcEtmLW9/3g8
E1CZQlal5llT5y/nKQczwoIxU+AR0bzndWqQxbP8FkxZYDXLgimM6WL1nbYq09LgOCLQC1R9TbBe
XAlzU/iz6Hl+Uhhxb3w5KZxP1BQLAsnvUubOwlsFkPVck6QpBCZlj4MFM4Fs6RdIxXWf8Mh15j1V
+1xGN3OcAsM724a17a3SkJLU1g/APYlhp9AMuHqFrFIdsYQhQJWas5E2M5VddO/2O92TvWpSMiQc
suHHQycCutXhDgUg5oz5iBG9MaV/++57xvnNT0ys47r8EsrLY2iZsj2wTYLiZp7NYr32y/QwZ9yp
OvMvmLB8sA4MxMSNwU8JGid69P9uJn2bfsBPVx/+XVaWAb5fsm8iCWhG3Gkp7ivFTn99o99fj7hX
G7wyt1LlBapdy7DbphLgT7PXhrqaXqurR6t1mSTfz23Nq0M1ZlbqgKguXxLg1zCBcrKtOMAeZo4Y
lBqSpa9olIoSmgXGl3LtEbJnJzrSXd23JYwX7XVvfUSEFRVJAYSiBVrH9fEFh7mVXwa1ZV0FwP+J
XG4AWT6h2dB3yKTjLgP+i+FHnpYQyzqkLUTtL8QqXDUyKJzPW3I9CbALtkJVaTFCUbl3HoVr2f7T
gqJXcdFwwkJgHuivo2NQsSBZSZUhxPeeMij6CBMQgzaKx9FYIslP3vZh1Yc/fZH80FJNuiERuWc+
QgPNt30IqBWE4LTiFVskbpiO37OkrUmMateMLbdrN+APK3lk1y3LeIsijKNI7GMLJJZ/ZtN2gfGj
YC9rkfCgjgTpdTTiRIxauOvNRqMGJfSjVUlLLOru43GW7/b2VRNPrZfXuVvXEXCj4kp8cxfwA+5m
oR1hj9N0kSNX/1HBFRSs343ET2DdpPUrPetBisMk//YXWo8mVfwByr4uS6la6D6jp+fFcBAMeUG3
nOmKRY27bSLzoK/RKmWqPZsPt1azhPiZQ//TwyJaESt1u/3ccHi28qFC7XxMNXQrricLX56br0AY
OlUqdoZo7919AF0xvc2QXvnE1ec2YTFhoVmjqSiVCHPI0XzxhyEKYj7Uq+KAQX+jvmpnvb6tkeJS
pjM9e1N2nBsMfUXK6yCfsOI5q84YqrGpwZc3fl/Rl/lrukPwCll/8/Eowb+ct8RzMyboB8UmFL5W
msm94oRBJsE9Vi6zKjs93R2AnEiQE0DmERqLTzYDCTAVwzrYDMWrgpWt12gPC79/VuySzS5+yUXs
5erg/GsiImdnyUe7KJ6K5WCvKKU+nGa2ZAjIbAQ2Br5QW8Ze8Std1N4M2w/9afJckOdjoLudBaiu
M1J44lqSzUrIqO/nB/nQfg86p6PGmHXCv1TSJK2AkYDv7I5f1nDoBcb/YVTGZZe0xpPqR72rSplQ
M1KFNW4zkplg8+IaMc/fpMBS5tG2kSl045ewSMFSrOq4h5VHNou0rDOtkJ+TldoI7TNmQy7qMufx
n4E4kC9+mfweIohq9oYpAZC8XRIYWSH1hkC4ovYih9ZWimdZoIoWBfOOiBfRoQila/BRHtvo0Gz/
sRRVFHrqe8TgPxU2aoYqxzxhuZ5K+1jdYcpA7XAuyQHA/tFtzNxBZh6Koi5LgmWivniCo1bqpv0V
7YDaGezVn3vSU7dVO6H7J2jDquUmHCFDE4Llu1CXZuLEGVH5OegBNkpm4dhxvottuyQle5osCsr8
AEYC5ucXzkddEm+qV9dHDh4Sg0UsUoLxp8aTuWi+lBCR4tEg0pYoNbyz47Tvsi1VnXW4UwCiWGX2
KUiUk5pli6Ty4EdNcJl/cDxn0X2Tm1b2AIZ89bpmgTWZVyEXteYPp1CW+U4Q7871QZW8kVIuBRCK
UGdC/51YUqdCG2DuEwOxLkbjHatoP4btNVZvW2FkTrcW+gZDoRMDEolTTL3KqvzVhE/NtB+4y4Xl
AKrovhRzhKLyqPTRa4nZZkpFq3FA7TfLUidxbTUlhCsvDKsmeT+G/dvcsIkoCWZExj14N9Rt8sEn
MDQV+N2XOC2y4S2nN1EadbHz++oxEGer2Bis6RqUG+JJCk6qCZhuHgWnTa1dAGl7z9Bx9fHsJuoK
FCbNSV59cil84Nkh9k75LTjfG8hcCfBtwsSatBTFJaya+gJaGbVoF5UgQkNWgM0ig4SiIIkjIj5M
gwMqM1L2/bpEPGLgJb9pxl15Ue91nQK3CPRzVbmM9LfPEfKpC8BFxzW5qtYh/kcSlJCpVfbB1vu5
IYeyicxeWlRpvLAgKqGEuzqBXZLv69tAVwkYQ6qVq0o76Ne15rm+fuyg5kqM34D7r6uzUZw5x6k6
Lu+XAeFIq4tKzwwPw7nsdXxyb6nQqfwD15utBvSuj8cRBZzZkY9YjfqXbGlA0fPbeYe8pGB6qBD7
NCd8vi7RVxBiOGfj6TNkd32NVROBwU2YV5FhzVpbT357i529r6Nx64OFAm7iuegjuxbE3sXIXeh/
8aauEORiRfrKAwhclGMsu+rl0DjFc17yzRAw5a4cScO0pK90/+mW1sO9AgrwdB2EfP/wJMSuv+gF
bZ91TmWxS3C0L6ely29urdkv84PB8r8bzhQN4UjZV/l67BYyfdggIqUXdHC6jeMyzRTLd987wVDw
mL+k0R7HblQNJ2bjByLVMj6thl+50CXN/qKecnEVE4qvrOsmD5I5lssdclb8P9HV8Kg3vCX0oSjS
V/3R3bt9zRw1Yz9NvwQaz2LJ93HtRa1ECGH/pw8UxXcLEQjRcc0YdDBOWfwDzhkkAPQ7iNpPPKKs
0gqiubeUCYLEDzfwCEgx7S1MMTZJkSnL1q56p/Xnpptw5INJn1FSb7ha9xO/pEFkK3hgukvQbmC6
XWTU1tQVXufDDSWmBAwOZNFHCSklQ1AJLMPNzGGAvc0yElHONToY2BozoekyJ8P5KW9dE6LU+ejp
fkuMCIxo26bsvp1S3PH9jF6r8VvSUNX2uAP7pnw+DCgi8D/KN2X5/XcgPqPnMcexbK26vi+4pyQo
9bYoecZyBOs0MouRgyycjN8AqUukwkJR7PQ9ZlW71wTcMzN30yX8aj/SCIWyR7LOhwwwQQCdPXR1
N28Zo2I4aRjE7gCK2u4gfgBIUmx4claI0rd+QtC7dBxlI3/8TQzccCMuqE6ippXvQ55AvOyG++SR
5J6QL9BK+f7YIgQsR92tsPLWco8vpizrD8iXtWaMBQm2bmbejluPTLOcFTmpmOPCdj4CI+cos+Qz
v9ypl+C1S7AvaiP3X/yVx6GOoQTk9N7AVQ6QPtVPfcY8ZsJFRFI6RP5B9ickm8X3Pm560Llm29KL
cEYqFkM2fQX15J47oaMMTtAAXhNbYcDW43jBLcJ79qSRVMcJ+3hPkWdLNZMU9c1Kphe+T3XTFV9P
uf4xnlmGepyysdgH8iuIDtOTkCNQa6txiBS0WZdcUeZ967oKU4mojc+H5yOFWZmUPG3gAXdsp9NC
welr7hIa3YBUXLkQWdIwijJeCj+RyZ3x8vYa7a9Rs8PYA8J2YFs72lWf80uDtSeC+HOR6jaX5UOH
q4cp33SBXRVIMIdn2DvbbcjbpkzpsYqTrDl6mF/V9dFHOG69QBQ2U27Qu8ayRwieKa65U6ci4WpU
kUCXQWPVOLjr05QG4D0Rj3Kf6UQ7TXEIFzvy3DZzzKTy8mCqNpvdgU73WdnGTFbSJarf4nbSUBJ1
boZBp4SeMlfAUakqidPSQG61k2179H3T1xvCA7uPjpFkjmx5GvSYLGelQi9c71o+vWr+m0dwWWcv
OeJxQfxIa/c1GAnMkuTb5jnuA8UYHiQeLd+UIuSF27TvRGdF2o9RxSOEnOFnGBhik+rcmxSEPrns
9UY54HTnbY+3nX+bwFYISBftWdAXymStlLvf7qdp8p9Q+RE+xIVrOFlGALu8ooO0NCHVoWS39LR/
9gAwGbHm8ywXWt0RyJ5Nh7FHs6EpdzF+Y1y/x9CEvtKJmLGqEdL/rCt8JWUSM8v8WpXqaL61Yb7l
9Z1TqsJtrZyQwBA1Gvy+qG2LzmIfoHaPn1Au2NttAk1C5f0D5WLEPqRY0vQ5wWj1AfXI5koH8EyY
Qff7jT+JcBKc4Ze6KztrCYWuzwbJE3lMWLdKk06nyD9hYAehcGuzpsBl2qX+fBao6cYL2s/o4yni
pa9DmX5SShO7ccrhE5aaTkKRqc2iV3bBzHacaNR0/bBraSRuxE1iZDJiC5PkQmfHIEir7fy8I9LE
lB7Fi4Iyhvo86U8ldDhUFTnTlnbGZukFiFP7IDp4rUAweYU8u4nE26tzYyIPWTf/r5wyqkaajr04
hS06VELr7klJbn41CFmGXVoYaN03Vz/u1Y/Xwj9t5MtudJymURCEssi6fAOp+Q9qRNJWEv2TQQ+y
ICTcEZX51KXyZbskY4MmovBQC3hw/ZFUYyOsJZbv0e+0ATMdHjBFPO05EyCeDNF8K+N97TLdX5o1
4foQmN3nyNQs5aQHXN9jJ1kgz0vcxhs7+XYAEnfl6DhhrU7xdul530Ga3YUPMKtrePDpTDncxnGu
slo2OwNWblX/JLLoOdI3jGM6ngueLz6PKIsk/G0GlFd18J0FZeMBVjmsopvY1xxwBboT/GcTReHn
VsMejVM+M96PoLUl75OIWLSAynFAgGZzdFrrqDX+gk/Qzh8EQ5CS0yMUJb1V0GWSf7PS3MVQhF5z
zbblhZ10zMkuINJvZm/6JFkSxvOlo5+9T805ERLq7wUOH5NdEsRTuj34J3ceelfGWDCVCmns9Wfg
gybKyNZroXiXD5Eoqqba+bO0x/Sp8C06dpU4UUV2+U6gV5xYtPndr9nJNsHU0r6qz+WVPLcFo8ch
NY4SFZpQ+tRERxTIBVMzTkoF069OXa8xwfBOU3sC+GCBAr6t2MgETnTUjGvJ5DCDSRXRXxNNfLos
Wo05w9L1avEfKVMIIIrax2SnOxwU4/zJrymfbLPG/HIpCEfMl4kAKrj4deUZKiCXSijA26GZQy4U
Yc7dzvokBjwDK8iikMtxNzekmdhHp22DEEgoIqLLjkJT7IXBjAHVuze12qYBOKlpUlxS4zNsmjwb
FaxmkwtxiTl15PCETF53shPqNjZEJMwTZCakq+gZmT3U++fEUQdqABO4oiIUhaO0L4+qN+J3UUvM
0D2kDpoTVHhA4h9J5dMyGxR778YdO7TSr32YVr1P1Qtn3bFBNJFvGJpFuF+oGBJKxecEkAJqBCoF
fOAqtYxzAb5VtD9x7NeEqzUQLYdtGBPvftFRVFDxfPa5ODkPRST9PcjfrbzJSSfb+kWU9XBZIcnk
5Ju5eEe+/zxW6Cwu+Vv6RCieeDaYgPQfxmjYig2IBvUwZ7/Ht4fmy2sDuvVKE3THUEOE/r+d1AEC
Y9+UttuPPOGqtDwuHJMD4/EhMQ2ER2Km0/M+s+cm59azNWh0CKLSEtnE0Og+MyryZz6NYnyoqcdb
zTDHKIAE7JNoJuLAHmWa6Wvt6i7J46hTcvfEwqMEasBPMsOJ5/aB7/L7Ei2EJpxujrWf4q27uEL8
d9O5ukdyBZnEIL4ERwDltbO/B8AA88CBaHml5exFpjgz7ULX1pkZbh/FYD7SDOFIIOJlUe0X5kf5
f9gZLSp5lgi/GT9XdypRLA1Qkh5TJ+ghRHGbH7mfkFvc+m0m6wNqz7s89cGgOGr2ZBm8ER7WrGt0
mPklbELG+GR+sg6spnQ7gmFYrRthugyNyOw067DvC+PjwhSDLko56utuzxrch7ERU3/RRYwDI/28
YuHMAm5YbmHu0mvKAOZ77tb5n0bU6qnliGwP/D2b6zFxx7vUkqEJl6Ynv3eZS52BQotL2fgZxdhv
INSYfwQTeYtmQs28QxxvnNCKzwONq/+QrVyO5M/+8tzs+6WTXj6lAhbRgiSkJSk/WCrDBaXu+b2x
X5ExTvOxkRRFohytVCNbzU/EIdD8RoXeILVQPkfD0Xa2hBURw3xYcXurCVGDf2WQDyuGdfx3Q5op
LMz32X/sAgud+9AghjTuTSLBxQzdHWWpTsnO3yNjEgx8h1of+D1OdB/SA/50jIRpuuP2XCNtPvjX
2v9bWX22f6iMzjTWuk3ruoCMXDboabWK7LSkS+3FQjWEWL2W56Ho+NQXmkd9QeL5m4Wyl24qteSM
Dfz9wsMxoPz+98GBwKJhA+1YksNI8hlBOLhiKR6xDHkVqz5Ai7heoCtAWZfoVDiU/HtbVoAC2bzt
h6dF6bZMpl9DwLJ5hnTjIK0jivv5YGAm6aT9h7nEZuFEDAa+DsPIPDlDzxWwjueHBz3c5oVV7VJT
VuhfLOhtCO8E8HfpExWgJ0xoF6GD25V4nhBTUhzLh0D6g4xTZ68C9kM/P8uf5t99OQVvVYVOCNV/
eRCexsWFUA8MGlC/51fGrNCZoFCr2mpx8DTYGIckPUB5p0OztdPLkHxn4XBXCnzp/a+ll/3/hyuu
VnY0FgmxAky58flfAXcXcVg0DC9bpaK9dDiIo8vM+1O9oHL5sNKkaCFI5ijiQtVV6LhSjQJVQbrJ
/8poPUU75q08ZnVF+YbjZ0LVDjMPWYCQ1D3gcG2uaUrqyMI59BKddenHs+lH0q0q59LTNcEGBYb6
ObvKooQC3pKFl1AwarU9n4z3ODqy7JqPFegeBa2x/4xCchC3tBvaJVxjX/anvqRmh9nwBkndwBHb
MTEqOlUbHIo1Eaj4xPrqiqRViw+wn7npAcrJbhWZa4fVodDr77BpCizzZLw5SuhcfMXHjUSNG0rK
OAW5X0tJzfjHMn8visxfcs551XPh5KpjjutldgwthI0gYfb1SdjieaxXIXGb5SsvdiFzbsFdgeBD
bN0eirjVMlFfPwBqWFZVp1msR61P/9KC/Dyay9AvPy48PUCp6CUBmSVWFjKcDDzAY/BSPKyx4oCJ
NnK1Frd6m7nnUV6sGUHOlg0KYXKf5mwyavzMJFqJOFuQVfMEIJX2toKw+q9fzHRZDoA4u3R2LyrV
xXmd5zFTsq2B84gbnpamCrFVg6NZAQjjZlo1OKA1nvaG0J2weUp2lMR9Ql0oKnPJNKhfZM1M3hif
Euh1iX6jmefVQ5w6IM9a4VKZRlq7AtuCANpxHACPbWtDO96HMDKv7fn9KswXTSF1bmMl1D4KJRfT
sXsrZYUhLjXNxi7EWI8iBl9tuAjeQa+gWl1gWpGrbOG4R/+JqaacfvgFSa3LFBW34ck0s+BAWBsS
/5jwlVE4mLmNjSKReLKKnj7oXo88DbWTsBOTEJtH+1y0dhikECwkBoZu30YjNtnVwL8+1+uQm4eH
Mn+oDqUy/KX+ZYO6Hsn9/1l9/tkmbt2iUSrxLfXMiUjj37BStixgU9AIjQGleMsUPHyNHldk0lCY
/8O90ruiWjFpJUUHdysxqhJs6d/cPcECQSnvk9XO8COHpOJMMuOEkzmOurIf8AXTFsXGJikZYhka
qJkyDu5UE0KXBm5hCoUDkP9/gCNKdrGIr2bNwQSyZYcqH9U+jvxgPMiQB3potFakqkwrF9LuGXo+
zRDRkwTyz7eF3DF9PB71J3KAqNG5xF6DbydtwIy9xrPT4UftLKzMkgYx2gQ+t02ui6n9CiCkhYSd
Pf33Z4pbUcZkocDJ5ywv5zfOgi53RJuNTQqD9e4PNjFSeN+iVXFr7wtYwXXB+mMEJ6+hWsVCGYe0
tIFrY58QQ1AsVq6NU8I3OE9qU6Fd2hGk0lVBexYX3gwAvb7j6tVd0SHmirw03/yvANBeAAT9xL/J
UMoSiDPmZcqvuEr2IaUtcWMkzB5mTHGuaAeag+C2q3HGiSg9084ENSko1VJylrZkj9ohsWmT8s5d
zdEH//ogl2GHVqMYV+WRNP7GTBbdpR6cfFV4Ua4JMV7z8TECWj0GkpMtjsdwC7tvMHw4zGrZm/Tx
Mu7O2QNshoKCaj1tc9nNfiPqwVvum0AlMdNbz//bVYnGwngHtkF3+5b/uaghn5Z6fKDyfiq0BX3n
YU3vr9g/Sf7UjRyzxH0zuN65CyWLnWravCLwt0DiarbRAHGvByw6Cp1FASxPXFIo2Zp/CmBz1B4J
6FcMwp2OVuXN9q1/2udIm9/1z6bS0IO9Zz3AtuPeuEOZl9oNyG7/1g9NLM20syoAi/ObygC8BE9E
EeeYG2yD7HkPmPL9Qbevro4MgAm5gpz/PmOH8QOx2mHkem9L1moR6rir5fQOjF85R1sQ1IQLBK2K
BrxAo7NyXKBA3lEWpEA+xwzTv3pwezpBFlwDmv9sXEiWWDGlvywXiGMdJhOD1m0O2597N8Q/M7+F
9GBt4d6vo4O7KAilPjn2WL8FSIGunuGF02rcz6dREuHv3rNvDzl7zqi7O8jOFwKM181fDT8m/K07
d7PL8d6aFor1su2lDOnnbgiD5UrkALRxGGQAd+AGROzMGfBVGJLGwMWfT2cr4deLlQr2hb/kKLv8
60ZjPsXDdGlVu8JPZ28BV7fMiFv7gmNmROP2LT3CK2pUrxcrA1eJsxaoASgWxDmpB4x29GMGYqou
TwWoc/T9CVKYTgv31n7X5P2djEtKCBx+BUeddYpGzYq0IyMoz6xkSaIpeNlXwNclHxoddqSUaTUe
jCX5TPq14JyjtGGoMQ1Z/vsLxbyrE5DWhuBy4cFHFAxZfPZlIfNqhLF2dLbiBE8EC34aPT+sXpf4
RlM3a8+S0R+v7qfqXW9iHf960dLwDTLnf5YkIFQmfxMpTg0m/g9EZea3ZR42BVffnT+zsxI2G1d1
5M+yXQxJVb25IaCl+Ff/fgsP/VQZYNB4zeiBbCqmW+3BjY243pk0d5B9t8Q5znqBJwqQLLFjTkxn
6TZON4W1u+Og6wxgHLxIELEZCrWCJ9NVUayVpB7JZvHC/QQZtkOVtRa61GnRyfQX6qzUDOln6AMz
2xnK3g+7Tm14WU2r6cdNbeVToHBmZKdhNZijF8A5TM8kq5sav1bJu/1l95XTO88O+g/wud/BoZ55
ZWk8FUaKSd2gj2iaumLlIK9/NBNsuuDEfHD+gnhW3+TCafyDxZx9tT7Xf6nIDDCzXiaAqlQFjbRj
QKJjRsQBxLmyzdq5CRvjRqJZ2r+ZZVov9+g9EiFDLhbsZdhmW/AOlY9pAbq0WH28g+XEJlJUuWsn
k2HgUW/oMoe9yzkY0vIOWiYPW1iKGCBMUGMQNS5szaD5Qp6e04fbceFpoOWnTIgqBY77+ezPhcLf
gwa5n8rorT0USrwBhS4PpCTCX/Mr/l67OH/zskvbZj9iWWEVRMlpbvAAawNEYr/rHRGLxj5BFCBg
iZoHrisqHk73iOCJZFr7u70gIghWTu5lke2MwcUtPCmUDmRpdUboMvlkqp/harIkfBZfAuBUMqkS
j4jvs2f1GISKNy+p2a/9MVqZ3lVZP3FZS0H2/pC3r2X6Lbi+2agWXKhusuFP8Jar7FZU/mWSS2F+
njfuMsbYPL+cNNBJGqWuLcf5RteGm0j/walwJaiDuaUVUVwXSSiiLRoOoCzjZmmhDLJmkvf7E/4d
LNZgO08R56sl+sgdpsgoi09y39UFdJNLLayVu1z92uVN9DueLwv3ce9rBb62czz3fwukBf6CK3vf
eW3H5xOTyTLVz/x0yfTu1weKQCLuEdqoxw4RRyepNzw/e7Pu6BFqNj189MU1fNJyo2qDAS2Cm/1C
e8xrnu18XkizHru5cbHSi43IlGQX1kPuT9B6LZY3byVZ+IlBc2e9X9nF3/EzIRJkEhlPuH5cFZoP
QXJBt5qQC7DM62N2tju7/Y1tNDTkmYhlId9leNQdydbUypuKHdLIj+j7ShtzvtHsgVGCH+44Cqpg
1XFNGSheukev0m4CsCAZuqv8HC68P9yKAFsIO9P4LciWmtFDdGuPLvbkZwZ+eqiBOZlR783OiYfm
8SSeI7O4bKhCWq85qlOhgfcbVSe9sFuK66bh557UIxsRoIx5hWa3H1FatNoaYvsO2Y11Ofh6H/BF
BY7stbqvYpDDSb5Y/JlovR5mSE3q8KGfGfwaKCem0R0VX8vB3nu8Wm+wwKS+HmSzpbIu6obKcnKP
86uwjZMfC7VdVDEcYNUet8pgtYg5Lz2zBuITI1w3t/YFUfbSF8K9Mk9UXs9eChPYSSZUlRIz6Rg7
28d08Et7+uGsiSCd9lO6sECLjX6dCQ5YV0+BpbjW8n+GURMC3oVXQaTvazJhLD1OLXPGhvNcdfL+
Vxb4HqgF/xQHL8CFiEhWrZQpstUnSKh4sgSyfVocIkb4IKIEp0EUI0U6d1JLVfciOfi3PTwCjUg9
C2TzBDymIMbfQXWieBhGpFHN0+3pznmwYbwvfJ1pfSImTJUXRExmYi9ChJh/G0dWlo79I9oVL34v
GLDIgX610dXJKyO+8SeSGvKnFbGFt+fOU1+HhrMDZdzINip3hEEcegvQVPf8n9JWuiXj5jvfNemM
do8lEsH65LvWxOga3ExTAQMDu9kBUYCqUtS8c4FJKfalomFcvY0WuCuZI82n16OKnHA5Ek3rKYFM
c+IehEOuZsxpGuBH2iU5ovFb/F288KJNCivoUDVBk057SfweD3KV+YskGicKFzYCNxb02sr7DYfA
Ehd2IF4nQTWhr0rJMxowh/YKug7FoDuClyo50sTYFB4MEjR0McH19QTLhnhG64qhhmMko8TG1bOs
txEZgWJDoMRit4e4bht6pi+ELAhyycINWJDJYpehSfNHh+hjG0GtYBCizT9wD30vEj08SzKh56Jd
5O/04LhbVwBt7WunoDFakCWy+0qH+WG9Gw9xXrOV9r8JzIYAzb5ciWl/WCQUtPfp3tGTM6R4Ua+g
mP+KSe2GsnGchKpuOcesjwClpdTnSost0b/O++3P3xbLpybPyup2gQeFPuzIrYWeoV9e0SojgbJO
rsWDwyDM2xwJAB2feJCDQ0ouWTKtfHAOjOOLOVmv9Ek4v1o7jZQk6vNHGd/wjZ79twwwDccqkpYl
zDNG73Fwl8W2mJuEAUBNcqQiXVNtF+SdYMIEK9duZRG2qehoP8QWQmNYBhYN5jyME4v6kBRruKLK
CM9wKbCzWShgri/DZg+MtQM/nhgXQ5Tr4XfISXJL6GKU+kik+obPpY9vMl92/KnZf0l5Aos9a5TE
6rWwjP+Zt2bE/NpGa3j7C1CjB9ZzvYvA2B9eqYigFMyYO6nxNS6h5gLGVXbKZB4vn2v9Ua6rQj6n
JPjqoO9A+A3ad5lwczOhdf3Vl5bmrLGfoGntSTuw/tpQuz7csalCKbpMl9PsSeol+53QQVpkVKfs
f7dW7v/YDtBCX2hkU3FDLqB56bTDamW2KhTulSIwRrSaw1zgmKK0gBCX8rrcJoEypJK2tqXA/D4R
vaLGk0HsGX4Z3gPycWl1GeZBjZnJnF8aU7IAZhnjGth9iLKVJ6Y1fTJlBN+v1/Mpa9Rtcf4fl3BZ
/yVDvSFHDaAiXk3W1QMyITW8Kkh2GM+RNihxte498j+pmuku2Nv1SIW7SpS4i/B9XjaSmiZyBnFo
C6McJmvLLGro7i5ookdokpFw72gAv2KHVA3UmuKOde6rxfjqtuSsc64QoF51aB8Ii38nmp8mLRAu
0brHeVmZ8ePgIu8BTGXMep8zx+OND5WgU0FGEWo2JYlPEBiPCGUThxshOSSpbEExIkerGXd5VCFE
kXQMfzLmveae+K0zshWVR94OA4mI6GA+yxYBF+eAMx98Hdq7q576pNIXdh4tMF0UOdnijceJxl/2
F38QZGZIKYOh52M0tAOMoVaGZgLQ0oK/hgmqpQphnDCnjrWO4ubsoiE41RK/sLz1MVRvaj8mUS+x
sFAkVVEv/iHzVy1gxt8u5bwo3XAu/Yrb/gIpEvCFhNrOjEatJ4k+ihnQVOAIaXaJMvm9aSGwHTNv
43/FitRly+/1qIVrRJIHk1G4ywvUDeXrGAV+xVLsoyO6bAn77fQlIv9Zn6MMiyVPw0I7atqgjuwl
NmmpgUXE1reZh1yOLtoVsF8pmMZMplHCw6ixdmoubQ1RS+ErtzzvsoDGnBMc31zllhs/xPqzGjYh
1PkKdQ7CZG8Yv3ifQxZdd9NjxETVFFgMiC9gPj+w4XGKs7nS4K8hGFjJwfEFJDmQa9zhegrB7QCv
WuluhbG/vnQRQqiRg8Yybzz7Ep9fd9uWxEyaDm/bhly7KS04SB9Wngt8ouBZxpbfyFmbvfFyP0ai
O0EPCVBpQzxEK4ohI6/qEMocfJi7I37cwWM+JyCrEkILAJbYf4bU8ND0Bf3sd8nUjZWoV1bUn5Y7
8zMblZ+GXnQdYfVbfspAS++hN2XayRmg3Yc+fzT63T9aM4P0UTEYn83PAu4gP2OiS2VTJWBL9gvG
UTOw6+TlxrrFY6Pb5NYrqdxTgfT7m/+WgUFXlcofCmHyQ6zyzUPrcqShOHS8CMVYwlstPN3TGLzq
pUAX4XbhQSFB3+mKP8QfrwrN26XYseeKgXEo40W7buL052SRylqEco7uwj1wVJEGiIJ4xkK33Grc
q+4iGsW8jPNuQ32rtGfrznfMjkcnDTul6ozcVTVPqar28VsMUay7Bg/w7nR/2NCQKg8HsJ/730gW
nQXoykOcFnPy1LijK3qPYRKFCuJ5DrDcxY8adJeTDkcQxWkloVj/T0gXl4Rgo4cEmRTKYv8Y6iHy
v2g9XrHTeiUUJXC318c3VVAdRKPaUxvP9ZdZerZ5GfmTjwGvHkpt812fc6TvuHMoF1pLhWiepv4q
eedGQFMDbVbNLpwGV1rUHbUXG31kfo9MXTCiimsazusti4nFXLzeiZUurCxOz3Lu7NfE8dzfcY1h
RmMFdOBMUZ9dMHH0/6KaPtRLYeNrri0YNyeWu6HrDITic/14J40uLeG3m2/ZfG8pgMk9wUWmwb9B
N2Z966Vld0d2K1SUYZEG98o3C0JaJLltfKvNFTpJY0u1WRaPjcp1qrqOWGVbTn2DpaEJMHTr1972
72E8I/L6LntCq9jW2nkQ8e02tetq1fjNfHTSpEGGTqSDof9wbwZq3cpxso1DcFNmKUTrBDYBACGM
sG58STw97/s7muJRCBzdG+JYs4DpZHetVcXCC2WdkDfxPhr3ZhNQBn5zSQg5XZP6h+PlFZuO31Kh
MY3I6YMvL6QViYQz7oDjCURIP5WORVG29MfZWzlhSsVee4PBdG32UhcWMDAN2hg52bAOkpnuroPf
y5CAR0+fTE/Bof7VfoV7hlztUOTZcCDUnlM5Q05Uh92+yDaeHD/vta446qk4EmtM9e/8tB6kjQ/9
JQvsp31NM0C0wzym3iSp+vmh5vaIKvaA6rSnhg8SYop7QgwugHWG2nmY9por1JYXD/J2ZiJ13M3Q
yAw8PCbHqzBIhiHwG7+Q+5ugRXnpLeNOW/loMCk9T39ILORE4v+3jVIWynqvWk7L3NZ5C8SxWoY7
H3lPlIYY8B9w2qTvYofbbwiof3HgIWYd7wKsLnJy6Hgu0TBp7QtvM+5m0zHgxwRL1Lh/lFAKQ8uG
wa3mTO5ybDd6L+LffA0Sd34OqtEAUeWDAK8Jhx19CIYEHRfe/4IBGydR6IRLDh4PAl9o769s97Tv
Bf0clb5bkUogqfZK2kEmAXG7aQ/SUD6xZzBOTK564ooz7jcXSqv167/B8p2JyS9CBCoA5NdQywEd
nn6IyMvOggDGebuGC9UjAuiVgawta8wuoahZWwjcNRAPziwH0FydJip9g8UutuIkDRXJ5LcvZ2Ml
txnkAG3b++Y79+BuhOoSGU2aPxXYZuRb0cXxxoQZ44xQuvFLl7dzT77RLAEg2N0kxXFDLOGG+VwN
P9FpU72Ez8a8CvwvCQVicYQMbpif809WNgrsrSkYaH69iauaKm9m4De3SMsbcIjPA/mMQzekwWHZ
wajcjnukZVLv9WSp0zee25zleJyKLo5Akq5w56o89uzHRdpge1v6LrjYSAklshm/LXB9lG7eIbcp
quGBU1zeT/NUegqQrjTLWUYJsYxDx56ysSX0MvevqQ3f1/I4GUdOUb8wOjInPupvm7yPr2HVGzP7
jEDJcSwg7VXP7mwO7loTHMNeL4SAW8seD1XTWTGdkWzjX6habF45/avu+gIsyHINZs3lZFAYfW0O
O+KZmeVTNUEKVMmNgod6mZVbeoeHMz9k1xHvX17ZFDv12LMa0nDdyl+Yw1iULl24yPvj5iAsV5F4
2M+93dviL/MhNWL0TDZ3OzieFpZ8kO1t1434cLyYC+gRtA==
`pragma protect end_protected
