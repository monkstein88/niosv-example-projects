��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2i�>�|�om�����x�]0�f���껞�3ւ��c��kc��A��|q���T����5۹���i8w�\[�ѿ��y9�o�儇pi�lu��Ĝ��)�Y\�+T�BB��-�5����֗�������ZƁ�� 6s}�w3�b�	�A�fD�Z>��r�Ob&�>2+�az���l�\�ܽJ� �U�pp�đ.8�֜B0���;���Z4�f�t�:?��׫��rX{A'"i��� ;a�W��%;�=��A��2(KW(�ܟ����5j۸��hH֪3I"���AS���g����A	����
#���oU��%�`5x�C��CD�e���9��z�ܵ��6[Rq�%��P�%���1;#s�2qA�D��Nޑ8?k��e�2�9n<o�^������i;���*d;�=I;�J?��3T�������Dڜ��k��.y+���>P��V��6� � Θp��!�P ����l�����1�BCQ4�v�9&&��y�!D�)?(��@���G����.�"�/��h�݋�Ϲ<3�lSE���סb��holٍ'�kS��?Ġ�_f��h���y���@ �7L�s�j���mB;=��S�v���x�\��;(�t�N�<��6\��5n_��#o��K�|C�}ח�F�F�Cg��/K80]���j��8���★������W��$B���W$ٖ�89�Jca����L}h��	8�@<�jb/��E�b��@��/2p'��V}����l/��֔���a�p�
��H�+�_���s�r;�D�l���|�wO��Ԉ��@xyٔ�6j�dD��j�R���$v^*�R��O�e�byi=�&/�L�$'�'����Z�|/q�F	V�Ze'��)�ߦ��}�(�"
4��C3\�Y����)/0ќ���BM�Su��K��cAl���3��>H�g���iT�gU��t`W��A� b���L4�č�U�^V\`�б6�K�8eux]%f�nQ�Z�n,�`z�`E���7cY���ɏ2@UV T^����ҩ����O��S���.k��%S;��M�!(�
���N6��4�m���'1����bxv�[�H���~��?�-sp,s��]Q�F�Tydya����ԏ�y���si�~�<�ȑ9����Ȃ��A�%o�R�����ĭ������f#���\��UuG
����$[��Ƀ��n��1y�<�>�g�9BX�+�O<�	}n
颾=+"{��ǄG�J�������V÷,`0���%��Qi�^ӵ3Kn@��!:{�4����6�AҒ�r*�����BRu�8�d��MHmn|��9Ka��:��ڹ�61o�`Cn,�ThMN=��f�9ɖC�̉��LDZ ��<s����F_M�������V�N&"�;�ٓ���HQ��Q轏!ݖrG� �����{��]��J3�=��T������aHG��̈́,B��1a�+O��R~+��)z����UB�4j<ߋ+�����,��Ҿ��uK=�㣯�m&�u�.�����֙K���
P�`J�n	��<��"�Ru�%�E���T[�d԰�����#�[�EŽ�Z3��n�o�9z���8(*�/g�O���ԫ�� ��tG��K ��aT�)��&q��6G��ր���3�%��Vi,j���Q'�賣�䑠��2�t�)��D��=�[' �!o\.��62�K��,+�x���}^�[���>��ޕ��	]6�C�u�W�ۗ����W0��C G\�y������M�T����z?��������_�U�zS˪և�ZI"dx6�����Y��� y�^�@�������Q�sU�Lx���H��<L�12�σ���bdV�\Tg��w�-Gs���nQ��L�k�
��)!�C%i�<K�T�FD4ή�z��8�ܔ�
���!��Y^/��éƸ0&��%I}�桞ݞ@+"7��֮�7W��]�ӱV*`AWEu�����эރF�Ί��JI��	�A͊\����	H4�O�i*O#�ܿ�Nd���0�WZISZ�<�')R@���;zW�h��I�E�j3��?D8xc2�KЪ��rfX)���jN�n�:����]��]��L6����#���AL(��t�^1FVp~���i�B�\W��;>��V�á\p��dme���+P�7���}h����c�{jD��ƽ ��SyЌ��[�����5��q�rݟ������|v�����1�~5�[E�+ҽ������҂ZM��sN`�|]T���q\K*�i}1���5�x�h9�*g�5��� �� ���u3_+M�����)�*O�B��K����/���/Bg�wk�+�L2�l���"�����$⪙i[�q���z2o�]��d(M��.	���u���Z�6�*�Cv�̆ݍ�����-e�J��f$6ۛ,���GZ����ߠ�fS���a?�K_ �K�762��-HPnx�5���jX,���y�͙!��J�κ��14<�o�Y3�y}o�X/Je�]�_ٚB�������f�o��P�j�Ӳxx`{���$��亢8<����tßml����6x�)�:���f~`�@؀�4����rf�s��{"3I��O�}�K��#��hŃ"�/��w�-��n�T�RMAnk.-�*my����f�D�]N;�n8l�7������%�9�ا�/��abo:�N�$L��@� Q�<�S��p���(�DQ��F1zX�j�� "�)��'�qn���$�7�G�v4]YFѝ�������SDE����b��|���C�̯�`��"y�e���`���/�Oʟ�1`u�]%�� hS ��@�88��Fc���Mw�b��ބN�	L8�;Tp}[C�ϡ��M���'�(Z��=h��*�@�>�p-�����$�"A��2�@!��H��&�1��s�f����Yߘ�4辝nk�X��<P �ܼ�$�6����	��g1��9���d��m��
�I��f=�;�\̑�5$�80����.4|_T�V���v���Yc�=�� ��V�~�)�����VA�p%�Q�hi%P����	���0��t��L�u���D��:�b�����wcy�S�U�z�w��(o�)�AZ�ɔ�a�OEbl�]�s-�@�zA��M􏵦�]4�NI�x"�:^��p3/�CwSS�=���)O�TM'ˤꊵ��^����v��
ac�^M�s��A=���;��I}{�\t?���4Ty�*�oMfA[+�����l�ж�v,��u3��)�l.�=Q^��`']8ӑs�b*-�֍�HZ]��^#_��۳/+t��=p���2�(��ɵ�a���ƻ[�C**���]��~ONG�I���p�Ap�X�����fA�17��DN�E�V̯��9��ƭ��� M[�����A��0��{3�QrOb�H[v7��x['�/�q�`�xD$f,�𚥈-j;� ^�� �EK�Ǆ<��=��L�tǳ3���֯<a�m�b��ZOSaƕq�e��y��CP���?gS&�_Q����"����\`�]�>`jnr���Q5��4�#�n%B���9@�|��w`#97踓.Ӱ-`�\ ���x@ӘP��8�
/�z��!�['�ș�!@����P@�\ �zl"����>^1�s!b�G,.���HŁ�Uj�W P,Ow��EAfHD��#�����_�oFU,S���m��cR�&@�Z��~��-VqaO�&D�}��S�g�`*�'�#\�	Kg�Q��=�����q��5����V���X~-�p��9ޯak߻
bz{��ԯ�1�N�E�Ԟ�	Q��|�G��$k���dU�/yUiƌ�&�
2�ymЬ&�l��[r��&0Nt�������*��%v�����R���ۇ����-�Fܐ똅q��:�h"O
����d5Y��u��sX���>G�QQ`%U�Q���/L����6b!F�g���ű�;@����K(�}x�E's�Bh���4>�C�:��%�w��:я��2Z=l�ͱ����E	�&Ѧ�fK����`�%����	�#���A�~t�����ɏ� 5����������F
z`+rѼ�zu9/�<=q����)pi_|&?}'^��e�Mh�?���#�c'g��"!�,�������4fvNϬ��/jzd�:�J&�ND��eƼ"���
��;��Pr��\������-?��d7�Z�Go��x5��D2����U�g��v�f�Cv?��]�O:��灀�*�3{�)��h|y���t4�X��ZNfX���V֓����`���������FY]T��)�r����X��5G

A���%���t�t���x��������1��hӺ �����{d�����	6���x"~�U	>����̐��s���3�W�N}ʳb6u����LP���F�6}T6]~�s�M��j�0����=�\��ɉ2�V�5�?F���q����8^'�����I��>�F�d�fim�y��;ۗ�y���mi�Z�3�hYC�v)+[�ܞv)3����:�NPH���c/�l��VB;p������ݨ��A�
(���B^h�P ,�el�
����i�|V���{�я��������^8��{�0��/����?\@��1)E�Q�� ��<���I��c����a�@u��&�?��@I��R�G��c[��0��Ds��t���T�B���I��P�$Ce-!�����|P��6�Յ�p��,=���o�k�W��%ȷF�B�Z�I���O<GX�8z՜Łˇ�(��=�FG�M��;���K�?�;d#Fq9\|��}�
��-R�������Ⱥ	*�Ɠ�Ev�y�F�݃u��m4�p�#��:�Ȍ�}Ky�T�M�$*0�����c@e.����9Yz�Lo�"opr�>˹2�OI�<����p�ҊJ�F�������G`�M?33��H��ٌ3�"w��7ߡrf��"���t�q+�%�q������>��6Pn�aF$Iw�����7��v�o|���3��Ů��>dt����1��b����v~;>�\}O!�/{�T���`{�|�s��+�װ���NxP:��1pg��W�O����C��a�tg��\јoQ �β�������B�԰�D߹��aH�U`L��g��ųh�>*iT�O�z��j;JΌ�o�;_�Nh���0��z�VG��E���42�9q��
��z:��n+�&c�@��͕�d��RF��*�-�����ͦntF*�G�A,���vlP�%��k�ޤU�^����?-��u�?�*C�{��ꑴr?�5!6���6~�	��KK�2q�bkJtH2!�R��Z,!�/,XQF���D3�?U�#���Ć��mh�/��d�V��*���v(��:���7��)}zи��Q��r%���e�5�
�y��4��[�h�>-�t�,ռ�g;Oh�"%��˿�[�pl��ӄ�l�gb����TɼM��@7��Ei���-�īV���r�.���`�$��ˆv�p9�2y�gc��_����͊�����WyPUt�v��� �DIz�������I�����w��!��%�,3
21mtNZ��C4(��M�,e�]wU�5L��.�^s���#Vg����A�C���*w��C��)�d�W�ry��DVd*��M��3��	dx^ �V����=c=o=�9���I<h^�-֮<���T���E�s���wF���"5G�z��~�F����F�W���D9����>�v�ahfw����`Q����d��8ۅ)�9��3�7´1�jR_ѡ�P8c팽8�������2�TӯUz�oHI��>b��PQ����o��L�UM�J�������M��Lm��3�z�4���A�.=%k�����ྪz�I��0"�s�h����La6��"�^Җ����F�9�����V����k��`i�Ōe�C�Z�[��Rt;0��H([u<�����N4 o���Ʀ���c6��o�˳֣,���3�Q5��Ӹ
*�u�_ËRO)��˵��7�g�k
�!G�贗�D��$����m.�?r��[�6�+�Yr�J����>�4f!�c��p�A܈���ĒJ!�SB�3R��zV��x�̲�$?d�Z���N��l�O(P�i��ts���Mܦp=m�Q���RUH���?�ٽ�N�]�K�F�����Wff��\A�1�8�Y����rej?��.�o�p�u_z�w�S6�YHғ;Q-;alU�s7)l���b��u6:b�-������qǀ><�K�i@��8U��it�>w<DD1�p�~�J�X�?�����b�+yBW&E��m"�ԙ�~�e�1W�?k�w�ղ��WU��lc�T�c�?,3.�R�-�x'��Ƣ�֕��+��}�J,v�0��O��� �dMa���ζ�Auo�Dj&S��Tß)׃f����.����S�q��O恹F0�� �;��Eӥ�{�v��wX��>�؞�ۏ���R|�^W���@潧�V<K�B����s�螛�V�7�鉘�&]kn;�w`ef�F}
�8[�%��5o�V�*s�XѤP�ѠU1�,Ŵ���� �~u˼��,|&�[�}�[F�-"�HY�"a~҉),BiU����<|0	�$N��eT���z
Fe�2(���1=[�K�B�C1Hl��ucu�)Mk�߆ t�NqM۞[�"as�;�o�>B6;'�$�L�zQTS�j�/����ͭ��d��	��n��^ϖ�
��cy���fihy��߾��3p����b6�������X�|X��U����P]���:06eq$wQI����/����NK�z��0���ޟw˳d�f���A�-�/�q�)��*_��`z`�-a�=�F-�K��377��}62�}bR�q�PSݽ;6����h�����Y�n����|�w=l3�&g�}�'���r���3��A��� Ɍx��`�|��&��Y+�/�H��?�E��a�����}���������w�<����Gr��H�$�(%׍�|S$����<x<b����:�W�җ����JT��_��4ʹ����t�Hr�}Y,��D�$$��|�H&�b�ҋSC��k%(DI1���\��L���� �v9�nL�\�H�-6O��x��mх-������[g:���`R�hQC�t�i���u��]\�r�ҎS�.�d��v�v�Wʰ�1K�ɗt*��z�YS(.�,����l�	��C��;ŌĊ�H|�vX�����l���$���͹-⃶����i����X: ���.B��g�vC�Z�G<�+�:5t%ޕ��Q�'�X���,���K(�3���th��?I_@�\�o]�/6^�!�#�T ���Y���	�W�{z�(@A��b�@mԧ��@��c
��_����פ�Xp,�77���`�g��R#4UI.J ��Y]�K�ڋ*�%�,���Ys"u��#�O%��[��n����zjd�����O1��z���Z�OXRx�O��G ������82D.�j��l�ED������%m��hz>2�B9�TU�9�9�1���$��L9F�\H3^ aR�@Z��M,�~�*�<��i����$1>�AV������3()d�C�OI�l�L+4��Y]�+�d[��?�\4r8��1k�$�%
�x�wS���Nb���Np�Ǘ/}a)�Wԃj3���TɮP]��Y�>��!G��>,f��uiUoT9�Y�a�5��{�pJ�VX3�+��Z��x��4A���Kn�-<��^�)�AZɅz`��n�?���CpI@�Q��BP�D�R=A�o9u�� #}@���[���9Ѳ�/���O>����֋=&��zw�H�\���~��I��Jr4E����EL�Xp�^5'J�t�eC�*��<b�G9���a?=~�Qd��2�UY�5`m��'��g�!>6ܔ���N��w�5Z�?E����V��e=������oi���N�2�RW�fK%k�-=�?��r`!�8�o�P�Y#I��g���<S1с�Y��(F8����,�!V`��X���N<�
����M�]7�K_�!��	bU��������������4��R4�ߌj$��m]O:]����E4<�"�/K���8z!5�H���JD�I$�i��S��£"91h���2�T�|�s<HN[§���^~{Yv�icf�膰��jm7�V��{�~��q�,��/�UM�����UZW;��Tmf#�R;j�2_`?qg1�"�̌}�NI�a>��(UR���jK/�ڨ�ۆ���FI�U�M=RF�޻ȩF�rxp���"�U-�j�p��k}�
��o~;�M�u��Wm�A�0��_�/�F!�x��6�*-a"p(3u�/�J�
h�W�ڽ�1sz�29�ʓJ�	��3qҽVC�`��3�̀��)�&��~�F;����l�����+� ��z`AU	4���ñ-+-"�.��w0.�] ?������Onv)7�xLr^��/L��M��r��zV7g?h���pY�ɳ���D��?$���f�JP6��y��s�:�Z���,z�:�ѮO��������s�2l�eg�0����K�PQ\~����!�z��IZd����I��eKE���.����Q�~+dw��"��^����Ձ�+]���1
Z��]a��fo o�<08t��Fx��L�2b��g^��j_�I��]�� �y�A�e�/�^�;@��A�W�[6�~D\��y4"����jFCC��f�	{�f��&.�Hxb]��;���"~��_np��	gw�V�\f���8�>w�k�*N��kR�����1VMv��8M��#:���l�>���U�f˪�my�\s����Ceր�w����?hG�R��'N:��7$�!�o�����<�!T)8�h!�:Z�O.�PD�>�u�\=Cw���`0�U������Fy޸��&6� ����4�$|!E �x�A��P���y�	#�)9D����ّ��وW�aS�X��}Di�}�S�8��(�IK���~P�
��ƌ������yڦ���%w��omQp���!�ẻ�@�B���+Ϩ죁���'���͋k���b%�����7����� 9�,A��%�m�L�4	�F]��mMԉ~ݽ��!@T��LȈ��̄��  .�@}A<h���ݥ�����2�bA��qr� ���Z��v���+���N���ż�߇YP�{��;*��N\�N�L�I�ש%I�x�� +#}�Ch6� !�+��Ee�=��_gF0��q�G4�}�u�vb���
��.�����&&4v<��o+�����1��RǗ 31`p��XeL_�,�K"8�\��C� K�p���2�6ӷ%"�ݠ/�\�;�$b�>6n*��*};�ve_��04�#Oo,7LJ:��<Mel����>ʰ���Y�Lk�U����L�<�"^C��9�(���LX�1~ԩ��MG�wэw�� �$ʱS�z��_'+44@8'���MY��O��q��v��R��ܲ-��E�!6;�l]��њ��`��ӸS��ߊ��������\ۏ5�	�C��'I'��=,��%}�#h�
��n��I��>A�c���f�n晰J�a-(�J6wfV9A^�۲û}<Ƒ�<3o�5���(7s?���ܧ���1@Xc�U����l3���ym�+ۑ�z�.���(��ތ����eʏ 5M�2�7�q��C��9�<��S��4�۱����F1����9���XQ{�,x@*:��ڰ�E��-���&������z5��.HD�	 �G��#��z'#4�Tsؿ[����b�XI.�>�%;���ؤ=:M�Z���qg�����u��jQ�. cb���x�hY�#g�5x?1腔ռ�~��۸Ιn�l&��nz1�=*g��y�+]����9_~`�Z�%W�!�ʯ¯Ø���@5�����"G`�|Br
B�f��PT'9�H0�l~9.�cԔ�_4UpS�+��b��}������Eu@ �Tz$�@����I&�jO���2�nBu�v�$+��jg�F6.3�_BQ�?!l{FiW�㸑�M:�q:��.#������c���a1�e.Kӣ9t�B�1~tB	4�]�F�R���
!z�Z}�w٭�I0پ㿿0ky�BA�V��7���<��Flb�*���JQ�b�o�+�t�b/�U�����ZL2�;���#��֡��{y�B�i4|Hfx��%���� ����w�}�p�D1�2�Fv%�)b�n��/���ʥ�k��ܟ��X�4��A�0��M����Ͷ���ƿ�ѷĪ2�t����q{籠����"�*X�F -���ϫK�@䎩���%��>��q���g�ɷ�����Z�ٵ*��;���2a#�����
�������U��jh]nFdd�`���+�/�M��n����2U�K��F�<	��{�I���F'��EFT���B�tOa;7�{��L
!��XS�MlF��z�7�hv�.{55��{瑱���J��m{���Y�W�νEl�1�u2�F�V��$7�m�K�A�8i^�mU��䡶0Z��fՔ"�}T��鄗���|��U�G�o����ĸǮ���e��U�E���ۗ�S�1�i�ܯ�OU���r�}y��mn~����;��4�=a�')I�=�J��ø�#������uGP&溆����S�l�e�|Lf�r���NS�397{�M�l���fi���X1�Xϻ�$��F��k�4g��@I�%�p:��ĸ 
i惄�������M���1,FFts1�9��=��p[���%�M 1x�9p7:7!�׭ֶ#�wWŧ��XG�!*K�M2Z�˳�N�O���֔��0E�p�"Z�F�*��S���Rlk:��dy���˸�}-F���`�{�aB��)pE�b> ������_aT.��A&D�A���a��a2�h*ܽOM�~H!��r/d}��
�1��>f���%��`T�~\W�����M��V�t�kY=2GC�&�Օ��mG����bb�ɲ��ZEZT3hMͳ�~ٮ�D�p��MR(w�iEJ*�Ve� T����9��$�ީ���Ea�Me,F��-�`���Dt�����Kf��P����j�2��Je\�M��a�}�i�}�w���C*�G�R:�J,�s�SX뻅׾����8v����7���2��=�͑b�m�'N�Ȩ��|��bNB=Н�����u4��v����!m1%6He��ѢT�!C�u�����a���#}{���kP[���BNR!б�����yc���O��H���Y"1O�p�%�3���)*\��u��X�zU��g�|��Jב3�"*��w��;w:F�[ʬ�$Ui��7�|Ƿ+=�3�!�����}ë,&@���F�P�ǰz�.w����l!��&+T��������7?��?�:6B���/e)) K�
���UX�F�P���8�UT��K�C'%p�Fm�k����,ioH��&ד�Vu��y0�3�5��x,xf�߹�`(�m��2Y	=}���֎n�2�'��hp&l#L4%1Zx��]�Ջd��ÃgȤ����s���Nlc[�eI��y.l$5#�Nj
#�/4�9�┟�1��4��m{�2([SQhE>o}��m����w�COO�x���>�}E��\�>B��ZҎvQ�,x[��`��)�����y��T������P#�*�ϼ�������+�mQ��ò����\��k���=�:o�>�8��ARܑRl��d�=$��}��K��7C�;,j�T��l����]�꺯�9j���$�W�D~-�]s��h�꟢�o5҂��1?b�_��Q<%�`���_�	�߫ZGA��
%���*/�)8p|�$Ϧ��|]0u45=��W�|e�`�O��4nW�&�l����3�����GLJx��>\/dep����3@[֤�K�o���� #JO�A�N8�X�Q��%Tҥ>��i���=s^-�8: @�]��ͅ�N�8iw�$���� ~�,�Q�7�h�z\���F������ck���I��}1�ӷ!)���!�g��c�yц�.��t��zJ��Z:Y1���db0���W��%�f��,$[T�]8�(��yǡ��S$̈����$j�[cNн�ĳfSS�ko����9G
��	YF��w���u*G7}�"�ZS�Δ���]�UG�KmϠnً;�\f^��C�0*䅀qV��C$̵>w|�Mv����j�p�/+�6,�#�~{�\���S�:_���8��T,�n�"ĠtY���\�u�}�c����_�	��!\�u���k�F��۠z]s(��_�����88��#��7PAqc�蔮bj�X��_H�k���PM��Ku&`���Pe�[3 ª�vJ��$�U�#г"\U��UG�b����,j3��-rJj#t:������-`;vV���&��`�f�m�=:j����S��H��2n���0�����!]E�k�	�W�lI�}wA��J70s�%� ��Y����5��}-�n�-UQ]�H�����,B���!8u�^�Q	E�~�����x�U(�����d䙋���&5�;�1�WКIW%������Ús�v�lC���['�{�@��k�$�R�G�7��O78f�.u���M��aQQo�2N �gF���Q
�S���	~"���z$��H��l�0���c�S���W�t���/1�G���=�pp�ɻ�<� ���ƪOyq��?�ׁ���5Sv�ݚ�Jii��m�nN둢� ���@n�$v?��m���¯�T�~�K`��1�������q�Z��sb*'�E�x�j���h���ް��@�KMz��Ҝ��\8Ԍg��?G����������ԡ�Q�_݇])�ZNPʡP�V	(~��l_Uos�$ts����QD�F�,�WT~�>�������օ����r��}�.6�,R�)���TRqjMPE���m���:����?jC'�
v�Z�>����Ue��1�	�Ɲ����_�nP4`L�6mggo������?�R]�`�C�Z����k~=s4��l�:��ؐ�e���0�j_��-��o���NE�K��n�@�}.)�U,e]i��*k�=�q�_JN%)���rx��w����eE�E��Sꕃ"V�/�Lͬ���aǺ�^�q9���#x��T�ǹۏ_S;��xi��@�>͵'��1�r t���}�J����(�!��9���i�O���yr���ݴ�Y-ri�O�/$����T�_ ��r��HbN6ї�%y�ۮt���0؈��Z~��/V�Y���;}�m5�`w�eD�j�\�?N���p�ͽ������vHTΏ������1
���tg�&��f; �ϵ����0O���D�g���;3�94�-�	���u7�|����_2B���c3���+�[oxX}S���)�[�0J�Q3�緷���UN#�?��O�zJk��Id2�����A�uS���NՉPJ�
������x��S}3ړCf:C�<�9�d��ԧ:FFo)�έ��t	�~�
;*��.��g��X��S~J�OG��k��P��������q�͑55C��E��������KsP;��r��T�J��篥�|��D�G�7�P�R/�8�X���d{���i�A1m�(���)G���9<�t;D�Ǽ�|�@"$O�#���l��8�ma����-Ѓ�D��.���P�a��۴[03�������x�������!h�_r�}�Jd:�i��d8E�C��Z*�E�d��O���1u;��"��π6b���LN����»X��[��׏��$4u&�Ǔ�D�R��K��C?.��V���X��؛i�����a��3`# �8`2�&炽�֮�d�j:�;��#�}�X�E'�F =�d�r�g'��� (�o*���XMm������Tx��U���FvfA��������[瘊2�t�P/�ی��R	���70O31�?��ģ\� |��V�u���gрA�ִ���_eTSx3σ�2#'bXX�pP�Z�г�����^!��i��z�����������~�O�?+/���1�&.��x޻��YY���[�����~v%yp��&�s�;A� �χ�Ѝ����p���W�zZ8>��]�4��.�����K�a[ugt������L+ _�C丅��6ᗲ�\�6�kh��Bv(T���3~9��1�L�w��JP�\��)������Q��i_y4/*<�Ӂ�����F�e��l�����dY��W�d�����D�:'wC��T�����M&ߒ@ܤoþ�<&j��ڡj��i;�~@j�&/0ɔf�w*g�E)4�	�d�Կ�PXQ��RKV���g*�F(����R|��'P��h���P3m��g|<�IG�luu=��2����Kp�}�Y��!J��r3�;���?%�2�ڈ���nWtٙ�I't[G��v��4(�� ����F���w�b�A�a(���8�ѳ'쾳S$h1r74-�@�.n���,���@:2�jYp:���b���{w�#���Z���Np�H_j+�m~,�fu�`}2�Z������usyx슯��r4`��8�p�^Q�I;�o��qbd��Z����G=�Po�U7v�N��%��Z@��JA�A�R�`���}�7ӗm٘�,SN�|�^�X+��S<fap�Q1'y�A���;�Cu�(��b�B^M��I!�>ʿ���z�����C�����pEDwq��?@S5���oo)�MG��I�n���`�(\������Z�	�\����eB�`4�RHk����i@ ���{��y���d�H�H{t�\M-����-п�?J�b3m��]��#Gh��9�))҉2��@R�n��i�W���ߣܓ������6Y;ZG�������&�;Ti��&� ���9�䇺��x[Ǻ~�c
>'[fG�J��Q���0E�9�Կ�8VJ����&�2�ώ]b;��J��;>ҵ����H*�O�l���"R�z}�u���x�q��S�=&������ +p���c�y���D��U�+�����;��P��0�<}:'���tO�?�<�nh�C��+U�_�mB��K��Y��9JJ�:S�q>ϲ=�5��������u�B��IOe�f~7b�!���$<'��6�v��.���XXQ��z����^�zF�9"^�K6�8M�F?;M,��_�����3~����	I���7A���U�E�$9n�t����]���`�b�A�Zl�3�IX��ۛy㍳�/5�U@��!�(0ew���Y>�g��)�n(����킩)���\�a	�!��*T�Ù6S��,��*��flԾǿ���= W�ɵ��:��Gȭ�j3j���"Tw�kb�p��;�2jsIe������1�!����;Fp���;�Gx7�s��%IL5��v��O�V�͆_Vg">%ܑ���xX����m��!Fl>�r!~�����=E����f�skO�d����-�5�<p�<F��4Ȅ#|���v�����lq��ʸ��]�ϩD�_
��j"ޟRbtl齏�Oh��2@L����n=2\�v�[�3B2�� ��2œ�q��~]�m��0��撳i��4o�;Ê��f~S�� �h3[Myc{!
G�>����� ��+��&d�JI���{���"�8�W >�/���R���|�\TB��D�iY�,D�l����񳅨��1jvxy��������w<�.b��d�k�"���k�1Lw�xd�h�!��A�����u琌+|�}���n&���е
��˞������(�B�TlaF6�=��`?�wm�:����99�^�m�g"⠉�?�
���VFcZ�P��;3�=fhs�_ID�I�ʽ;����`E��.��&��C���9���=���h���x}D9Q�G����6�S�.����?�����3��Ȓ�����Nv)8^�1J�����u��X�� �� ��~VA}G���4��}���:���6vP
#������{��W�2�1�^�*6��ܓ%�&̣P���b/"���j����!gQ�?�9D	4w��֜����R�a	��lr�S�e>C�q�������M��/]���P���Vwg�DA��d��ee4�nɓd��-��-;�x+t�^��p�:B��U�����c�֛%��e;B�Î�N� E�7�<���W�٬݃7��8˥%n�T4�4�o֥��=��M���2ĭ�#��F;s7����Ŭe� G��c%���Ix~E��P��	%�{��DI?�*���4PH��H����E�NOs��Jx�e���>e)�	X�*Y�j������~aA[��6��&��-t�o+
���OE��_����$]��ŃEuW�w>�D�	�P�\�L����씡�%93\��u]����>��UN���Y���@D>��u$"���j�v�uS���1b"6��������>5��	;������Ce�-u���W��n��L�����џ�eg�w��l_;?+{��4���h�Q�e�q@wַ�pmE���䏢V!�Y�����_��xh�f��i8�ى�#pI��!Yql|�>?��k���&�K�B���R�x�i�ܨ��F�����)ݝ���i#��ϵXf�TѶB����&�bl7$q|�Z��i7�\���"=������$�b����
�	nNN��<h�԰?f�'x��I��o��b-%juPW6g��K��]8���)�S2�,v�k�ӊ�ʨ,I�u����xŢ�BR<@-8:�QDa���>j�ǆ�1�{�7���u0��֑d�q}?��Eu�R4�h��`L�J4,�8���0�?^-��@��QU�7�V1�6
M��6Ff�&[���2�04����70�ˋ�iw�io�0a2d}C��o7l"]Ù ��Ln��>|��(��-����5�i0y��G�=q>��qK��k ��@�u�UU7�qu��V��'W}O`��m���z�����%�Ӵ�t�/K+ނ9ٓ%������׈.�Ṙ�$ӥ	Q�^9�Y�3T��R��O,�k�K�⸀���X��J]%�ڼ��p5�������p��N�Y
!�-�&h�l2��9�ۙsٜ2�\N]����:瑤w��mӻ�|ʀZ�U0;;%!C� ��4G$\��h�_�����O�Mʼ����\D��xV��q��P��I5M�V�}��ʸ�NO������z�CK]ӍI�j��$Cb��R�2��ޓ��#9e7�َ����2����k�Eobt���7�R�;F��H;K$�Y��2򦺍�siON~½��p2s�%ԫ8���
m�jY=�=KI)�ȯ��\����elAl�T+.V�?I��J)l�L'�F��t�T~N�w�v�!�,[�M�
(:���n[�^��#=���RJi �6aR���5��c��X
5�P�(�{NlЛ��I@��?���9;f����\��%-��:m�",-� F�w�X5�ތb�eWwi���͓ݧjWam�I7F�21���\�ռ���5h-��1�S��i�*�YAv�*�H4,>V�.=Wy8�c[��$�
��脡{^�t���S�^���\����T>��M�L'�cgq��O� ���d�r�"�l���I��u�M~A(¬N�8�~{����砩�X�?�����1q.��L��?�*[��=#�ċ��Ī�h��t�?+�pc��k�B�zDA�GjTA��X4�4/�����cw�S��gێ�RXC���(�&ֶ��i��x�s���=;a�17Y�����Y^���m��n��P�j��KÅ:�e����SӉ���6��]�'g���4��:o��s���wb)���?��V�9bI��٣����L���5��;���쀢V��S���Ѧ��G�T�:�5���"�jFUO,8eL0A�,v�X�}Uʜ"��pQ�3;^`*ϤTmڍSq�c<{,[h�!6��\R�T�H����I3�n1
�ؘS�r�R����V�����d�U(6����`�<h�3a����~
h��Y�\	]QG�L�':HyݕG�C�B)k��o���x�	m�iu������O̲�`6���4`k؆(�1[�?�߈�
sQݷ<V�u��i�LptGn������/�o�ߣ��N�/S�q��ּ[
������	�̕A����m�H�T���'C}=�0�E�U���ʹ��}�ڬ�.��CR����t�91���uS��<�0��c�*t٥�q��DL� ���CUG0p��V��R��0��W[y6��'~3��|?�j�������T:�Q�D���^�}��y��A L5�O�S�\��h��i�����'��٫�xB��W�M�����\�6|���y�g�:"ڟ�I�:�0/�TYGW�w�����￳�[�!�[0X@~5�<3�ZQ�I ��ݰ�8
r�8xF���+�[�厣e�g�G����w �>�gR�¢�zL���Ac!J>�I��'zT�]�F{���Q!WץƄ$0�\5rKs�����5��Qp��Ӡ%>��6�>KC=�4
���i�M��m�>i+U�� �B��ܚ��^=�|�f(��=�^�`ђV�e	zet���L���F�.wU�d�"1����(��8�O����+h��hG��V�f���8SO�T������ rZ�{p����ސ��y�pL���ʳ�U���4Q$F���=ބ'��$B��}fމ�dk!ʤ����1j[����P�9$��.|�r���9�Ⱀgۮ�\>lbo��s����� (�Q�4�x�@�����ǶHM:�z��Ѵ%2w���|���6`��	's_�'"��
���ތ�-���A)��ʾ��
�Eσ|'#J"�V��!��X�Y_7{�y��)����*�d���+��W�q�"�3ށo���`g�E�nQG�2��ـԔv�<G�ә5�S$���3Q}O%X\����y��*4t'�Q���p�~r�~�G+�{�~5m:��A�=�N�%� ����!��~�_�)ç7��v�wi������c�A�kA�ԊR���|H�E<��?zSa��]Mڌ���Q�ܑM5�1ؑ 0�#&�x
eQй�^ �7҈]eh���S�)��F`.����C�"d6�b�>�{AD�~kc{�C�1�r�m�5�8����L9AC��,1[��np�s}n��T��;]%��iB�����/���`���=	 �i��KlP-)�<SA4\��Z A@)=z�Ƞi��I����71���k`j�>����D � �U����g3C8�"�	!kD��y*���p������d�2���� X�˺%]�u��,:ގ�[�i�V�v����b-dٕ9�����P��1�l�P�b�W��!�CX~��iK��ⳝA����<AYW*TNe�x_����� �.$���B�Ǻt2�d,�V��w�C���[�w�ו;�"����~qUw�"�/���.�r"�l��kN��d#�{dV��fUHl���,4���69��M��v;��B{q�Qw��(�.q�GS�T�F�	f�=�\����h�(�.�fǧ/Hf?`ٲ���q�pe����?��@�g�+�V�3�LR��U}�����1��0�{��j���9���sΏ�1�Ȟ�<�c�8�8Z�pU�FI��2k��m�"����}JѽKn��C����/H���c4(U�)U���1�YS�4=hX~[d��� E05����3L�m�@��]��t��%mg�@*�k\��'�-����J�l�,�E��}��R��Q����{���&)@\�ES���0�h�N���BGȵ�sH��f�]�F
� �[l�����3wĢSaas�����5'BUVJ�#/@����r�V`��.�$�ʠ}ϬW�]n�:Cr�c�([`t�x٣)���
�.�6̭��7�hq�ՖBX*�T�Y���2���5�M��:��}5�0c���]Q�+���B��D`J�����AJ���ϑuE{\h~���g�8#�1'�3�v��h�jHA��e��EJ��Ș�I!:|I���ƶ�"���ʪ7��b�|z|�n�lq��]����ۤbv���� ��Hӹ�`*����3u�޾�I�χ���]Ix�����r i�P��=�2�U� +�y.>���nYˑ��Pe0B�S��eYB�r��i!J�%�f`�THs�>0_��fmV)#]2��"
�	ÅJqcI�T��֣�8����<{:7?}V�g�@��UP����l��d��U�/o_�������!Зj�0Ɂgb�'f�;5�RfX0B#����#u����
(�E�`T�Z�|�"�d�p�7]��J4'�j���/��-u����5]9u9JLѿ\��_T�����y��J�����\H���>���#(p0�(��l�͌!ܱ�?m�P9�&����/�K)�j:��_�0z��e��i}.��-^Ѩ/S��Y*ȰOb(�o&���iėPv���2�*ˉrvp�ecU=���e����w�[�v�xΞ�8p�/M�b�	C(ej�-�0sQ�T��y'K�WwnE�%��!������)��U홨o��v�x�O�8>�d���ꁚ�Q̌�kˉ,����H�ZU`�˂4k��K���C��Y;�?�8G"�:�����KFy��,�\#>X��w��ّI-Cjl��_�#k�B���DJ�;�й:Xᶎ�̱�A�쪎�|�'�i�̶�9���u�)�v��h��k�Nl�b�kJ�q7F��!�u|��l ���Tf�T{��������(�xp��G�(N��ԓ���+��Fq�����Ui"�C�w�0�� 
t.�Y�����^���2G�զd�Z�D��0��[;mv�C��4s1���;-�Ɂ�|�7�j#��݂�b*�c����|/&��&~�։�8�z_�?���
��U�k2R���A���72�J�҉Fj�p/�<��[7�wШn�u����A ]��4�ѣ/e��U�6�_����f��uB��Y�g����<�.�mR�:�M
�G�I�e�ә���_aC>N�odD��?���|?\Ғ���Z@�1��v�;��ĎH�άٞqU=�?�ۘަі�!��(]�'&�ߵ�:`��}f��`�ӝ��q>�c~h����z��g�|{@�Z��G�m�J���t�V4`j�!�d��D��L��$o��/%�K>lqQk�yJ��^݃Xz%;+�<*����e0]j>tr�˼�����|l�K�h7<�0�zI�v�?c��n5O#x�И`�Ef�T}���{�#�h�IpIw�R����}ZF������yPe��dz���CF$�۴ #!�K*� �Epl�|'S�ˡ�����0ל�mb_U�9gy���&�y�S~�"�|�|R���ך�*�vVQ�Q���»N�$�%��L����A���D _}N*�#�!S`���S��ݿ�`k�zP�l2NThw�D!�&�tR��vKK� �l�rߟ�n2#!�?%&g��Ѳ2?)�hҬ��Z�vr]�&/1R%�� ΀����D���}K�x�I�Jl{�� �y��P��"j��_~�z��-\��6T�,��"ٲ�����͈�������WhFw�f�<�NkZ-��:rԏ~�5S_TF�JU���=n�A�O�R���/
�o�פG��YN�}��*�^b��mx�+�|��\��W;[�)8�y�宝?A*t�1��:��wY�D����[i��./ـ�ӎ�?}�৞}�������������"�c���1`�}���
#��6F�����;��A��u[L�	1>�����b��<z��d����������C��[h�	ՙ�UK���j�+ �Ň��+\e ��g�\4�P݃k
�Z�l�%���\F���.�^=I2
�I���w��ck:pY4�b��K:�Z�bL�c���fD�#�$���),Ճ� ��?�љ�+6 !�S�
¾o:���/G�-Ի�i"�]��{�.�H�S h�T�޴*p)K�z��'!�G3�W�/�Q$$� �BY.LR�$����?���Wa�e��,�y٤o����z�]�8��RZ����K��y��g���6����ڳLO!@?A�@.I�"�|�7���늭q���+��O6�fƷ�ڷ'�W
E�i۟/3�sx���U.Vz�������ٛ�o_���`�} �%߇�G���\�DF�輬��ܕU��5i§0H�q�Җ�D%�y�̔S.���r��q��z&_|¬��v ��4iDJZg9cS�!��}[i#��Y�m�	��LH�j��3e�5ڢ!rf���t���*��Q�ˋL�1��1B�G�sՏ�.�u��u�6@\����$<��Dm,�ɀ��Bj���!�#(dm+:�Si��c&�֮��B.O���o���+��)M�=�5�~$u�5;BG�����5�����6s��ں���,'�B�?5o�n[���	'���2�	��N&��5��Q�^\ϗ��em�'=�T&b~LX�aJj6;�)��^+��D1�{�pڑ���X��[�ձ��u���x��J�M:�����x�5��a�h�5F�ؠ?О彐	�	;�E�#X�9��c_��UM���)T�>�&2�LX�ц6t��Y`/;���u����-�)M�Z�:�ǚ������c�Q<���Ԗ�/ǜ�>��I	n�Ê��Sq�<�����xz<@�C�e���<��-�*w�x \��<O)�s;6�y��>h�$OZu���s�Pn�Z��D�ؤx���5>�{��s�H��C�u߄>��A>�Ap5��l@��$�~��CY%�;�V�4i�.��n����B���ean�ܿ`��^�H�4����{�8\Ǌ���W�Ӛؤ�_�;����r? �W����f��I2�������0BL%��^"��#����D!kI	ᾓ@��e_aI�Up��.�ZVaZ���8E~)9#�MhL�Fr�������@#�)��R�J�[:Hu&r쌅�WzvT=A�&
9��7����>,R����3Ֆ���z�E$�)*4�29�Cg'�Kg�`��d�*,s`ɪ
!ј㒟���l��9����3&��#�3��|��o��?��u�7�&bP����i��P��C�\�@F}��=��c�@��h[�"� �ĉOW��Z��;�]O����dhn�A��a��!��ͺ�v��K1�!�'�ͩ�ʆW) ҹ�k�+�>�)	Q~Lڐ��I�W8F]ݩv��a�&K�����ߧ��A=�T��û���N�?(�t쫥�/F�OUe���σV���C~�?��H�;��h�v=�V ��X�U��a�3d����MV�ó�
��̸��Ѩ!kA^5���T<�.K�aF���,y�a��� L��
JdFgD�-s�<}GN��O��`�RY�ৱ���-6B�l6�B]��B7�m��q�+H�I�r�m�Ö����ż�cZ�WY#�T�r����f��Jf��}Yx�CN ��b�C����E�S`G�wb�Ti�s�+0�I�z�Zp�1�PI)h��]^��tO�S	�|Y�H����,q�,�.��|�SMX)�Z�Q�;	%��tѩp0�1��_�KY��v��S�=ئ&w9e�3[w`4�ݪ7ASi�Ӣ�T��V}pʵ��Ͳ@\s��6G]���@!���Gڨtڥ�B��k���=�#*��n�����8�Q����D%}� �qk����������[����2�������9c� ��5�sqi�m��zL�$+��hG(Y&��6=�X�6 ΂+�{����E�$ߞyp=�Rbha�sJ��磷��龇�ͳ�|q�[Ř�C���H���*A��pb~ˤ��HO��D��ͳ9�o��#��2�g�J0M?ϽI���휣���AG/���!y����3h�M_0�k:�[$��^���G@4��w�]�_[ @��.5�"�8��{�!I����:GG��;��L�3�5���f���N���X�+	�`kPH���W"q�<6��|~w(P%����4�������*�j!
���-�N�cRRhx�P�D���nw��+�~C>��s��G|A
hm'U(�MX$4�UbCh�����EZO�3��M*���a���Gk��*���+�.�����
�w��UcZ�V�|!2g~� �i���8�K۳ii�t�5"}��4�hd�
'�g^"F���7�����ˡ���ðG��R��x'�URv�;�4�r$�~�ړ�s��To�h2$�=��-�dE[!�D���� �Tsg�4�Bf ����ʅ9%���N��O!M���	�;��#���������6{T!����t��XD�"�J�Z�4 4U�Y�c����a}�Gq�7�qE|��t��޴�b/�u}�K�V��-F�B.Md:�7��������N��'�x^s}���q���x����G^��\A0蓨���4	2���	Ȕ,]��\Z���-�r�&���n"b�8�~���W�_p���{�� �r���g+���NC�o�?��brsLD�9�����^�� j��Q�+M}LUc�`�e������|-�fĞ�e"�Gx[���s>��*�1������'���>���1zŐEC�V��K e���å2D�<kϊnv�&2��/��p���s�Ȭ*<ޗ��_\�)�F(�����hbPË����Ջ]�+4�I�#nz�`}aw|�k̎=J�n��}7)�f��m�Z�\�s�ӼN)^�2c�2���I���^nJ,���H"� L��.V�h*��KV����a9>҅ۧ�� 1^��0k��~ѓS��d�r�?[�T�Y�ǚ6���K,fq��
YT�L���ִ����Z�WAH\��eFM�٫���y0��RJ��	��j�@<X3	�f`�æ%��� �@?~��l���ʒ�&����t}Y��fb���>�I�|i@��%��!f;ȖN7�8���M@b�ι�
W�]a/Ɗ��2���ǒo�Tl��\-
�Oњd�_�����������Dƽ.�M}B�9ܦ���i��5<I��k��j��ٳΦ||%���&�9R
u�����@{]˂��醃2�l��P�h0�����p�����m%a��dsrl"C逦��ѥ�\�w��\��F�bͽ��ϵ
��L���pD����k��i�b�#�l�lWS�#v%�4F���6��س�|9�ƝW��=sy����W	d�:"��1)b���~��$G�	7{*D�cqK���*�\q����yaY�5ni�@�F��l�������Ga]C��9��	ʱ�_U4���r����(1�qEϡ�_rk_��	�J4��1m0W�$��IX��,zX�lϮ�gE����v���`nH!
��S�q����[���8g������р��H��R��u I���c����i�kޓ��H=Jg'��}܌���qon��Y�I䂬�`�~[����Ŀo�)
��K ��-5�\P�VJ:�/���;-,���iz�8����7����B�0�K^c)�)�`V�5��2j9}[��>N��!���'�����m�F��^��\��G�2����nF���i�c6LCb���*$��;�3���#Kp���V\�������5o���?�����x��߮��mQD���v�>ΟO)�F�f����pF
��C���˛j���r���ғ���x�ܚ\�H��g��l%������/����6FRQ"NI͇}�@ۘȚ>:��s�fc�BT,��4ԹՀ�v�����(�PO,���fD�J�o��M��l/��ZL?A���0&R|�w̣��-A�;�\�9ԺᘟGFL
[5c�%r5�SE�|�P��cmg-�+�C�!8�
�w|��H_߷���J�+�d�������uN(�'z��5z��/7`˭f�����B~���Ǩѣ�-�������	4��<�g2��tG`��8�+��k~�.Gbj��
��m�ܜ��sｆ� e�^���pH�gVw>�j����z�rZv��o�p���ۇ��y�=��e�7q�ά*ǳm\�๒�+�(�+��Y"�����sc��L�h����X��0"^�<�7�=ص�v����m��^�}:��O���м�ฉ8�	�%O���Yt�;�إQ;�(�B۝����;a�_����P��T-vX�Ȉ�v��:�E�lk��
b|7֍��!M.�-�*EVB��!�d�N��}aTx� ���Ǻ�^e^fՌ]e�]���i�����(�yEŸ���NZ)���%���y�]�������.j��(�ß��KbC�DGۧ�s�8�f�.f�=��Q��唂5��>���E:���ć�"<���u��l���)�;;-pG�����s]	�g�#	,~U�U��n���{%� ��x��r����C�Rq����Ãq��F0*��zR�jd�!�����X0���^��K�������6�C]9fJ���6OQ(W!�?��|��/P0�����b���Ѧ��/-^�a��%�a�ܘK0Nwj��l�߻T��IȜ��2�+W�7�2��u��MMC��xS�퓥��#%O���d�L�[��t�J$(}@x�H�/
��!�K�S���=�;t9'->i�Zk�j+� �#�S���1�)S�躤�kM������l�Y@�ʗ���:$�<�����3m��l���,Le��J;$Z��o���l�݅p:�2۹'2�/��+��n3���hVz�n44����d��ϜQ~����cB@_�����N +�s�k�_��Dј�)��<����z�~�J?���~P�n�n��#	�7����ф�9��mz
F�Z�n�u��"ؚ9ȿiw�çlm�'M���g�(���\Pf�1U��Ւ&@�/��/��x���Q$hh�Y�F,���CM=\�Xz��f\��)���c�����XC����W���=To�ߒG�'�������=���"|�����:���@qnp>o# ���ho�%���YPz9�j��M $��x=�p��5�Mu�Q��<�Qz�> �rU���������u��&�Kn�i';�oLc��_��5e���}�?##9Z�o'�"��S�.�}̚�0��'��D�2F�D��D���لs�c�B#�^�^�J��4��F��OH��%fŦ�'$/)e9Ä�g��)JK�/n� ��t�g�K��6b�&�&����nn%��휂�#�e�ڢ��m��r� \�g,9�S`��KJ��7{F,'�-�z�S1A����Ud�` ͟-���xj��0���6���z7�>�ۇM����	��E���P͹+F�t��КuQ��
�5�k,Ds�+����E����r��p������FV�Ȯ��,�K�vޏ�~ĢD�0`�]L��XB�u�a��`���|N�a����*u����A�q�4�=�����$	i�*�F��Y_+w��M=��M5s�S6��[�dBn5u�^4��T�C��`�G���S���.�Y	R���G�n� �ܟ��C�@�s7�|��""�X�O;��_�~$���,�U�q�|J*�nm���$�%�* ���|��2*��F%4���C�Wd��S���D�;�������xLQb���8D���gq��[���f�l�ˆ����G����Yt�dT���,zX=��T�c��hn	'YuS��) L���Γ4��7\1��7G%�?����E��TGs�����S�+Bw�&�g=�uT��
H:-�K��;�x�jS���������ډ�Y�Cc0#n�=<��N�//5�k������8i�Q��M��B֒#��y	WD���,7�M��3���WF��n�,+�K���	a�E��Q��J�@�W�$ї=�D���_ �8����0���`������e��(J�������IB�K)��1�M��a1A(���W���G�T�-Y͹M2o��X3���e+�C:O�u�,[yǊc�{��?�UV[��Zj��l1�@
�ѯd��͕*tD�4m���Y�9ە>�,Ü0��w�Њ1�4cϕ�L-WD��<�1�hn�6�c��'�)Ox\J63$��J"/�G@��{V�����W�oI�#�N�1(*� ^�H�=�4Z6������N�zw�<%DK��`�)U�l���
� ��L�9��g+�e�=�����,e�rR�t��XyC|�K��j�n���	o��~�;�g!�	�V׼�=� �e��`�������\͏FU�^�y���B�z��^�[Kw,I���-��"��:�傿���)���M\-����2�3�fg�T�|��C��d}�_��mԊ�"�[21D�>y��G^�N�_/�Q������*� _����H��8�[�&v��T��q)�O+ه��"=��i�<��C�,��7�� |�>T����O�������q�m�#���H ������Yb���W?�°����fW;�F��ˎ7m����ouEU|F�iSQ���o�Cv��R��ct<�!�5yB��YDu�Gh}4Ю���(du8e2�`E����~�I����V-ذ$vB	@�F���1�BH �	-]�~Z��iRC�Bk��X�T  ��[bwu���on:V�;n�#u�_���޸'�NP�ߔ��`��Y6�D��y�������[��T��ő��B{���'�^����,�_�xo��ۜ�Л�R"�x���MlX�azF,l��)E (=�vk�`5vG�-R�U*��\�=W�`;t���]��}|-?�t|4YD�+8%��Urxt_7���~|���ߕ�U��p� ���	k]�Q��]�����I�U�G�[��?�hG�x��B���!`�[s�,"3�q�0M�S�o��k�Tg}����U��v�/Q��1n#���%����z��`/������Gb(���2Y�'�'�������2�W��g%�&�n�}q��Ǟ��x3��� R4k�1"̵�R,>�~�&'϶jMZ����N�}r�e�ӷ6�_�aeT�_Iߗm�_�w�,ET���S�"�}��h�S�����я�d�X�X���1"���Ѵ�dŞ�h~�� �C_n��c��o��wYT�x}�Qq!N�;ͺsE�)V��mʘ���ЬM� Y��ǻ&
;,Vf.־[�4�V���ض[>D6_��\=.a<�c���-Z��}����<�f��ä�W=���$�Z�`�(���q���}o�yL�sU"���+.�P}@c8���"m�'����SF���c�!l���`�����#�3���5x�C�ο=�����a���sj�_��݉�2b�=��A}��v)�!d�U0��y�epU��?�r8~����V��ӛ�b]*SaN�Ҁ*<�EPhČg���H���G�EYa�$�{T�^�V�R�g�y�5Xm��g�����Z�����c�����m;��P4j��h�DO�qa[��|8�I����l4Bc�.k�E \SO��'��!�xP���f��D5��<���
�b�Cj���P3�I���Y��$j)E�֭J����u���38tp��� ��''�:��~���� �=�������L�� ���=%}��ӇU4�i"�y��a��6}ر�:r".��>F�J�v�<�ᢱ�}��Z �@&4�5���9	Z�����8�0�ކ��2�Qzw��/M&bX���)�O�e0�ZN�yC>���;H"^�6N4:��0	��& %m��v����� ����3#��j�E�2��;���׈ٙlh�=e3�,���<��рé&ET��T��`p����	n�7R��׍��2s#���6�W�k��L�z�D�k��z�8�kc��RO���/�eX�����Y�3T���_8�Q��j[l����z��������"��n�ˉ�G e��O�N���n�R�G�\-�����h�K	�K�i%�X$ԖI�ZO!�fؽ�m)�Ii�4��x��������m��~ws�h��ح��U�hqqx��i��y=N��k�f�	�`�������5U����1TF���!���h�$�j��,�9�m���������7�B2�Z:���WUj���U!��Γɐ��uӳ�����˃ty�pB|����ж%�bl�� ox�s�f~h.�^ơ�d-��YN)j����25:�g���p�כⲯe��-6)U�Bmd�S���O�N$����*�9M�Z6�^�LS�5�8����Ӆ�c͐yFd�t�,��AƤH��P����rBO�:�����Lϼ�h�,U9*��5���JͲ�mߜU��'}���P���I)������[E<Y�<��l�H���ġ��{��{x����8��}��1�ߺ�B�����F����Z)x)4^�#���oL�n��]�,3��;#��m V�e��O<M�>��m��T�W0Aj�#�εA�Ќp"�3��n5^P���g�~8Y��a�m ��l�SS�� ���0��^�~0�0<��g���3��Z�)k]"&p�9S^�¯X��$�U��d�Y� !���o�$L���\9��/o|�h������R%� n�H=v�l\�	M�VL�&��Fe�Q��I}һu�����=�ʽ<���b�4/�e88������b�b��'S��LT���I��ȍ��w���i�#��d�[�e5rh��ɊS�k�����Pg;ryl$X,_�~�� ��|��7W���E�����tD�V�ZB��Q���C��e�]@���㧪��R-`Z3U*X�ȑu_"�q��9��xN[I�,D�'/�Ő�}VE�, ��d��3���a8��o�<^ߔP2�V֪�m9^��w��]|�d/�I>X�n��ShiZ I�U -{
4�q �8�K �����2~d:�^�Ě����+�T�:�'�f�vL��K^��??��t6�� W�����_��
xJ�pԞ4l��P��9w6B��R(5�3����V�8�BPO�C��I��`p>ԓ�b~u�?7�O��1��~S���4���0@�s�9�EyX�P=��.6k�)Im�en��d<��*,zp�����Vk�,ț�G��b��Eq�����o�?%��J���n�*��ʔ��������<��D�cz��ݏ����8�r��g!���Q�W;�9�b*>(s5a��sdM�$�Wֺ&u++ç�IQ�B�"a��W��͟�s,9�	�,�+9�J�.q�U�d��@���5�EM����34�l_�o�����ꑝc��Xf��H����#��ц�U�~��,�X�$n��TQ��
0�J2r�zwXpׁ�P�v8�z37���'��p�M�DO �"��#��I�2-���y�O�w����8Yg?���ߟk�W]D��P7�́�_���PQ]�GU=<��d����!�S�@�qI[���JG�L[��nŒZ�O������
j92|���(Ld��)��'z��&������6�,Q�ïKn�[2F�Vw7N�5U�����~�yLw&o0���6�yǣ�A�hXR��
�L0�iT��9[�!�/��g\ H��
�Ìؗ.(&�u#Y�a:D���&��E���Xͻ۞̡�Td�!ds���:���Ut�IFۿ�ׄZ��!t_R�o�W�F�-پ�|.�����]���d��������~\}���GB�}��گ���H��g��ê���x���)F���,C?�01����7$��9� ;���w~s��B 6y񈵉��O)f��.��^����"5xv20������\ayō�nS���̺<PusŖ�3B����s�Y�x 3FŬ1�t��U�?��@� OV�\PG�pte��a�j�����Ϡc���ָ�9�e�#ĉ�JŲ��E���L>A�	�x~P�) �*N$����rN���#�X�z��]:���^ǅ
i[s�A8�#�V�g%A'j ���^e�Z�MH�i *�&o˒�<}y:�5|�Hy�S6穾N��ё�).��Ȗ�I�ǆ�~&}�,�/w��i�)���P�F�7����Q_ռ*��_���>�iu-Y�MY�\���Ϗ��2_ �\�s�,0��:�Qf;��[l~�Pk�����f������zz�7�h�4]�Z�|ɓ�2d�
�=L�\GD_�Ϩ�+L���l������MKtM�,��1������i�E��qb龂g�H[&�;��0m�l�l���6��p�#E�i$2��յf��p@���G'�`�iN��������3C�L�� Y��/�/�y������_n��t6�4��BjC�{�B�O	�ԗ����!�itr�#��}e#���yF��b��Vz?�Q7��%ozt0���F=�����3�!g!'X4lTW` l(�|VV��		��Fs��-�Ʊj&��ԪyF�9لf�)TiL��x<~�q(�P};o+��+�Tj<D
9)��as����q�7E���نH�
��� ��<��yG��D|HR�� ��3-��c���\�� zj���Pf&5�qmٸ��ajH�i�b��h��k|%�;u~��G�2��D�^I:K�Gj�C�2����G�'��~�����/�!�����f;a�_�J���%VV��5�Q�o�� ����:��$l�}�w��V�jI1�N����x��DR�����i�l�qe8g�+a�+d�p0G�H� ������� �*��#F��+l�$p
VF��X ,�nx����ͅ��d���Q��*��yUU����Cc*��=��������.*��x9;(���<0el���t��v����	�1���?��8G	��L�0(/E�_�"Yv�W۵h}�g���F,ճ��x�H�pvE��8l!J?g���O���!��L�|�� e?%��ké���ݿ��O���&��.��-�	Ƕ0���E��w��]�e\�b��y��*�J�X�Z�l�3.q�~������������c.8�`
��*|���Ow���Ձ�r`�G�4u��y~��G�PR���;BR���e�J��K8��׊9/�>w1"�`ۜ�8Lwv�+N�}'��(y���7�0{��ŝ0��Xv�
�,�J��*�{��#���&�t��Rb�y��o�}\����c�ۃh��U�/����M~U�}$�I!�q�,bĞ��'-��[�^���k��sk6�,n����ʫ��!{���+h���,:��!��3���=�-"��ڕly�p�������r��Ȳ~]m'鳮H9������� �O3��(-��	����D◳r!��P��ш����as�	w:�P�R!����b�cw��V@m���D�ƕ�K�!�+�t�j{���p�D��	0�5/`Z#=T*�Q��ӥ��ۅo��D��|I��s�%�*�c�aG_�rͫ�>l�B_C�Q�)W��w�a�t�QR�)9!X��Z���t��覢��T�ݟ i~��)��uoy8^�;��<MSJ��aÁ���ޜ핞��+S�`TF6J�����N�����M�4�F�8���ͩ�8�<WN��-�o��så�R��?Jı��>�N��I��v��f�nBn��t�2�� >0`���c7ȡ)و���<�М«<�� ���6�������*�3���@=\Z�Űzw���c�.��ӑD������!4H�gR-e)������O�*�RN�:���3��hZ��iC���>ه~�I���s2aP���q����xZ�]�4�Jԫ/�5�Cał����0y�t�.%����qt��	���H0���[)"����+�>!>�#dX�E0��:��Si�E�J"hyt =�T��E��,��"��jÅ���yYn�6�W��Ԍ^BAd���4�ÞR�����*��tj�n�&�B��R
��^z�}�V��P�[&�O�-�0gh��ٔT�	<cB൬��ڵA`� #�3c��Ǵ����[Y����h��A@��3�Ĳ��51;��+�>#m�s��Ǡs�`T1���+2H �~SC���:C��Ɠ�ɚ�Yt4���̛6@j5��U�]{C���T�c��ʩ���p1
��R�O�8��PfW��ËV�h��4��<ɀ���/�C�L|h��~Ҋ�h
���cC���7�C���>P�Ԋ�R�%�IYf�'�z�LuH�+����\��d�+�ʢՎ�#mQn�J]x�X����}G'_ț��=�ʟ^A��ޭ�D'�t�\�֡���U6$|/NT�U�Qm%���)��ff�4�9�`����C?8����$��꩑�ڣC[�(t�����0�t���]�l��rvP/P�]����ﱹ�`eN`����I;v�A�{�]����wo������x��D�_��)�L����1��y���ƿN[��o��s]yqn@#�b
���1�#�Dݹ�mU�_�&~�=_:�΂���f�u�f]��_ꘉ?O&�5��VW��H����!�H��G+��g�T�2���:�} P�H%�p'"�<���N>�s>��?h5��mp��@�3� �92�J�-�/$�B2��&�5��o��Nk���4��YAj�Ă3L/K�i����l��S��^��:�$��I`8���b���Rg��l�9�#8'�XC���i�rQa������2҄��I�Z7�]�F|���<ƾ�X�S}�0A�?y�-�J�; ��<�{���M�G�Q�e�-{7+����/����Vճ[}Ũ�p�Z�R��b%�)E�Y{?��/��&4�.^h��'���Y_��x��X"ivt�z�%��]�c�t_��o]"~�%��L*���A�+�-V��y�eFA\�3�P1ءo���xѺ;'H:^�nW���v:�$9��R��'zk�pŕ��u?NSg�P ,$�������.)&�g ̹�)s�3k,��x���� ?�ћA��QS��Z���p�����X7QQ��l%6�_����������D"QÝqق����ğ�l���=�?�I��uSi~ffi4/M�K:qn�X��q�`��F>�>�L�.NR�:��>:Vˁ>.�RN�^6
qc�-p&����p;l�L�ȩ`����C�gƢT�m.4��.�埍|�I�=�AS��r�k���vA�Z^��)Mu[]����N��v�o+I�e{ջ�9����PR(�o�`�M�|������

a��ڝt4ZIխ"\PRTyapT٣��6��oľCA�_�s)xC�N.x���U�����e'&T�!:�7��5�ِka@�ҹ��8$�ln�ɬ�)�����UU|�(�O��V��T.���.5Z�/wZ.'�����Lc��_�O�W��_�>������%�.Y�����>��>{���0��^�A��U�BGr(ܸ2���w �3�砬�u����a^s6�6���8����^_;�,�X���4}]�+���
�i�]Nui��Ը���z���X�o����7���,��qߍ���.��d��N�0̋�QG(zW��g@��#&cW����z¿��g"��E0��*��b*���k��A<JuaHٹ*�S��n��`�`�,��v�_g��p�F�t��K�4_e.:^`@�xwI����̂�9q��8�ԯ��#��2���n��E����T|n�!���V`�3z]Wm?b��Xa��M70�"�Ml��_6��CBk����	����g�k�Y�mP�,����0�t*�lc>�7�uz�B�s4�DP�nͫ^��ų�Q��~q7�"m>�GHJN��KYZ�O�1��]��pg�ݪ�o!5 p+;��p����X0G�t����W��2{�!�G#�S-��Źͦ6"�@�"su�4�ݲh^�烄��5��U�ȃ�;�tB(�ׯ�͇Î�k�TOj�s\I��8#,����2IЊ�m���#D1�Iʈ�P���,^��ґ���Z�c�`��d
���u� |�w8�z��>� �K4|�R++^��*Ǳ]I��<(�d�z�`V�����3@ �L���0\�-�5�f�"�������g���.N����Dob�.��f��8y�d���	>��5��?�Q�G�y���/����g�I�
����w�`�3�c�X<g�@%%�ə�+|�Cz;P�?�X���7�3��ڋぺJ�B��o��}t�}0}��!����#3{�g.e㬘4�xr��.�MZt��F͌�s�=�$��']9��5Z��s҇D�g�.BP}��	<��F/�E2:�Փ�|��l�=�i�٘P�=��+�SL ��/x�?N��e�eç��f���B9$l��}�}��_�Q͹sğg=o����(��ԏ�`���%�`���1T���ĝ����R�/�pvٛ�Ӓ��4�a���>���ez�1��6H�����Tg�E�\Ús��U&[[y�_8[�se��4	��!��U��'�*�3�P5�9T��N�^lN��ש��[�U�-|�V��)@C��JM\|�N�]T�D��Q���� JJ:F�>A%�f�b7w�v5��%����Ǽ��B]gv��0����u0�@b���E��x\��,���7�bC��m$����Xdz3�����6�E��(�9�e���]@B�����U�ы�]��hPkB��T�,��xs��֌͕��{�sp��Wـ#nB�{������a��S8�?l�z~��IT�Ur�����lr�98���g��eyN�u�bQ&ڞ�� �?���g ���!=������*��~���Y^��o��ңϱFOO���:�{�w7		kC���5�7��p�=����d�G�4�qsx�c�)gR�|������t���d��������է!bp�Dq�_5����h���_)�Դ|+�����cDx��F޵��`��_"���_�
P,�o�rǴ�~���ׁ�d���On�G��Z�b�o� Mb�<��ء���9:��TtJKGC� �O�G�������<�csq�������<�8z�/Y:�%F�ե=A<	�P��t��R	����S'n�#��ɉ.D�VJ$��oG�[)K��v.S���LO4���m?��,8��&[� �K��J�3D`[�[�<0K��~� Xuz���M��#����8�,@��茛T���9���{��]ٖ�hy�ĘjD�ӷ�ul�lgH��:�V�"�^A���7r�f@�����Y���,���f�|&��5�\S��K6��_$�����Z���Xu�8Q1Jk�����.��q'Z������M�V�C�}Y�Κ���.����L���JV�fZ*��'�L+���xˆt"
���5��a��<��2&�&}|�[��97�=8GF�p�?��4��Fр(�`É���w�Z�(�p�Hk�c�#��k��OYjx�rURu�aAtI�H�R�~Zg<��f�i5\����+Mҗ�k�o��q�q�9J�����T�F/k8����?�o]��I���i�d�j�!O���:#�J�4*�o&g�㴵���B�w�ߤw̴�.PגB������䰻��%�G 迿'��6�(��/����f����,��^���s�J��vܪ��h���b�0Κ��h�
IO1���e��8���} ��P�1
7�6�|�u�33 i.?[ҟ�^�&����ng��RMj�Z���~d�t�Ό��T�.SR��Zьh��e ^�ɻpn�R.ר�Y@����~W�Vq�1�/wFq�o+ �⦕ف�c�ȵ���5Ш��VP��9о�aV�U �W�e,1��7:����	�T#��8_���HLgLvz &�(1�ʂ��)q̉ǥ���j;Rˣ���� �?��%b��}��)|���8�AX{��2����	sY�5?�R{ו���#�pV�K���ق'] ��|ptZK��Xjeu�PJa@X`�R���_���tI�c�a	��oi���J�9�@�c\4��ߐo©��ջ�rE��#���H	��t3�T�E�e�H��ƹ����$n9�>��f�E!D5^ߡo�1g���6A�к�󜉂T�f�Mo���:���M0#8� ��`n1�[m��)dL����������uh�x�������"d�[ymhn�ѭ�5��~Hg���5��c��}�ɫb�T\�v_���(��vf�k�`�V?��� o����w���ErEg�����iJ
Ah6Gx�J�u�9)~���QԺף�%��{�4��a:��k �Lm�� �Ih��� �ZX~���ܔ���*�p�9}�>(�}���(+塝`��x�����Q]��S��8�P����B�V�ȹ[����_�����/�B�\�s��oP|�lH<MTm����H�4ck�}�<���vk�u��x���-o�B��~/�LD���c)��ܙ�'��]�'C� �]�_%93��4l�dWV�xF�>o�@!s����l�5Y���x�x�ZG�͎a�&=�ϲm��2�7k���J���L���c_Y�u*g�y����X�g��w�5x�d����<ȥ/7�ތ��Z{M\މ+ةC!��9�b��Fb��P���1B��g-	:֖q"<���.q�`��o���?<NRx�NHF"eVT�R�.��#O�1����&ȟ��9�A�;b��*�p=4�ѐ�2:8MORfazY��`\,S��T�i��8@9�ޫ�{��f�ˋ�@{ۺ6Y^�Ѩ���9Z>̄6�Aľ�f~�.w��/E7-e�;���U��_�?�3���D�lg"I���N���gz�3�A3]�.H�&�_
�\()�܀���۩/G?8�/go�';V�W��w*�jvD���;�X�+
/�K��2�����JN���+��Ė�<�i �@��Ǐ�Je��?	�'�
/9x���x�˼HE�nZ����݈�Ē�� �mͯ��E��M�d��n"D�������yz���R��05aMDP~u���e��a���5�¡�����A+*�/��qkŘ�(�9~߀(_���"�5a�C��t�ff��V��YW{F2�y7W�U�廞��;���qH�A����՗E�9<�>щ�Zk��h`�٘0<���P�'�Qb����	%FY�=���L���s���>�T^Q��w��9�&9�A���|��aBGB7��I��Q|���:#�1�,ř/J݆��	���'���_~?JxZ� ����h�[�L��$VE���c����D;�j`��h�#W�I�C/7�>+/5y[n&Bv��. �3�҅u�*���ǵaߍQP�ހ��:8�#���=Ƭ�<�2�m[R�̏?��WxҎ�{e���q��i��������A�������'������(&^@�0_�u�CK^��BbUZ�1ߣYHZ������1Nr��b:��y����H�n�2;�
u[�Nޭ��i{��G�O���kE`j</�q�sztW�p��Z�6�������&�b��@��I�*8�8�G��_E�f4��j�%e �M;���aV�7n��x�i�a���w��f��@���f��D��L�'����$n(�|�����V`B:9��~�/�k�,��".�>�e�՛M��lt���w�=���X�s��z�Df`j�4����d�u�r_/I��Ip�$�뭔+NUĦ3+����9mS-ڱ�#��]� |^��d�. �?���I�r� ̯�����4�z�n-��2��{�X5�:���խ#�i�@����C��{s�(��>���qo[��?j��z�ک��BX|�E�-�2�ߏ��]�8J˺Y���>*��+F����B�~�V��LB=,���L=? T�2�J�0������n��O��9]O"?$��Y�h��'_��&b����SC�OE
V A{S�_�nw\�"RQ29a�p��޶���5�w�j2%f=:����];����<8��S����]�������3X�':0�ZSג�M螏����⛬'��g�'ΡQ;v������%��~��2in!�=y���Ʒ��W�@&�f��|�8�̝G�.o6s��5��<�|���ik^pv��*m��-W����b?p�y���D�\�J��#�T�G�dC���1y��m�E���t�Ȏ�s�nz����"�OL��a��Aݨ�,�߬I����?j[%�uG���t���rY�:��"Zm�g�T�J]��b���vJ7���~H�≪���I�P�̈́���du��H@&Lͬ7M"+WwHz�)cH���=�����1`���ДHa��Ԏo������$R�pE&:��Gy�h�h�+*31�����D�����+�l��񎡪�����=�ܓ�h�������2J^Ng�ťB)��c�l�95:J�\Kp~�����<�z�w���^ʕ���4xf
�K�4f+���L���X�����������a玾��'��,x�I�)����,޾�s���t���!e�_��u�������韨r��%�,�G{���J^Q$��Xuލ��H=��O�D��6hFܴ�s��3.b���r]��@j:U��Y��n'�9� �3X�v�ɷ�۰'I{�U�f)��	ҙQ�5PW�^	��GJ,;���ѫ����"Ԛ$��Np&U�ƤT�*���3��+fb:0��7�����}�1���A6�/�ܾu_0Q����+�Q��͵�[�L��h
^$�s�����K����Х%��alx��N3@m��Ms����aaQ���.���X����l���������g��&�P]y�r�����(��ɪ����j�&�h��ʧ�����,sZ�T����h)�(Ȩx�[�Β=���m��&�0�\>!Mɡ�x��y����]�~(��x$��@��{�2��x���N�f�X���iS��L.����b�\))M�
��+��V��a�؍��D+d3
u�@�-><+d��͋i*n|:��1� x���E��,���9�z5%��MT���
:	��a�o0{��J@U-?'�U��_�e��cP=���+=��2	��������[Y�(��N%b�p���y�F`70���v�^:��(�h��@¸�����K�P���K�oq��l
%�_	G($��4R%ۤ���V1���~D��
9�VYX�S�&�(5��9����}�.6�Tݚ��A�B��J�i�:���/��ks�����V��=�!Z�CZ�1:0�I�����ș,�('@O*����6"����<0( ��f����.Y�><(�VؒoP9�a�>i�p���C���u|��>m�Xh�c^�ѵ��u�@�t��<�';�C�6�����CȀ�7�"�� �A5����Fj�<"҅�P���K=�P;�*5�K,\{�W���q}\�#kd:դP3^�IEBC��-�����t^��?b��dUrQ��x	�̺��6f`D��	a������9�Ӂ��Saa�\z��m�3�g~�τ����X��|�w��+�������gu`Lq������/wU���S��xa
4R=>Qz����ͮ!D��\s����X��<����˹	F����j��f�r��,�N.�Z��wA�,�-h��[�i�����x��0f�����c�y ����'�+ 9w��ڙ�QS��8�N�U�'ȏ�P��?u�g��X#N��,����	U.-0�_O�i	�CD]AT����Q!�Y��G��$\�򮙻`!�>s���'�VܬN��S��/� ���p�͵�܉hhе]�awj��QNݑ:t-�/j/E^��w�������֊ҌX�OH2�=�k��ItLǋ��#�}�����p�X�ɉ���n��Y�[U�O�&��b�4�,�c-��#/��$D��	>���]�ſ�8�7��Eϰ�&���t.u��e�s/)?��O����tA�=�W$C6���U��FV�Z�w�C���ݳo �����fh[���>�C�tC�G�?��v�A�[�X�[��:�$FB�"�i��<cam�3�s�]|Q������Y��w���%у�;��}_�,�r���>9)��ԅ�9�@.g�y`�O��t�Ml���h_2HA�������n7s�Mò�6hB&jƮ�PkYA���Ív2�>�/N!���mS>�zdW)&юb��1x˵�L� �ED�-x���"jL��CiI�E�=o�%8���/�D\��8�O���`U/'u�86vL��9w���O_7�cG5h��V�՝�:H�E���c�GR!��V���YpM>��@�_�
��/c F���[Z�~�t$�d��è�OnO(_{���)_���u=�9���쨊�q����:�7����?���M������Ɋ+�e��3�x��D��I��k5d>�a��>J���~õ�ￚ�DM��򳫅v*)��4��_�
Yx8>�G��M#�J�c�ZvU��<�.`�t7��Ք-I�O���"����w�֜�NuɝUEW<I�i�%�#�~9���4�3��6���#�)b_5ڵi^圴�OҌ�Ѝ-cMy�a�`HAY�D��48�9����.,�
��Ǉ�y"��t���u�JM�[��S4�i���h�_/X�ܷ�k�|]8;Jc����n���F����v+�3ܖײm��l3��6��[M��)Yd��XWb���ˇ�$������c���SpX�Ϩ�CzBi������{ڝ��b���	�:��O+�`�'����3ukp�>���C@{�����u	�����/�]a�,���)G錯U{W>b�J�S��y:크,�5�_�/�[��e���IH�6���Q}����pC�I���tZ��ω���@�1�cЏ���~���a���C.���v���(?.ffl�r!��^��eU���[��O�xT��VԚP,I���S�|Iy���>���#��F4}c]l���������SlP������J�?z�\8� B��nd�,��J(ʢ24��kāC�6-�����ׂB,lv�1u;Ə?���+ו�~�p�<� �)N3Il���c�~�wCw��3�	��϶p�v���٨�x��Y�J��ݔ����a+}��3>w��L��miEO4�e����XJ�"}qs~�t����:��Q�c��y����G�+헅���Y��"~(��f�7�SΊ�C�5���
Ǝ��m���+{�ȣ��7�+�I�oh��q�9�,F�m�{��}]k��T��Ff����XWn� 0�?$j�Dv=\o�-idi=��q[�6Щ\$��M���^-�T��6:c0��>Wv Ƿ�~b����"&Г��ᑚ<M�]��"����҆�qMW�(	7��a��i�@4�c9[$��.�7�U�p�a��"htΛ����%���i��u�.�zU��g=�3�6fW��?�B��Б��%y��z��'v�Қ�t��OIJ6\ !��x��*��cVp��������k᧬�y�~O�`���\�D��y�8؍p�@H���A�x=Tu�e����n���G�>�|���*�f�xE\�.�ŢDQo����eoP�$N@���TEijV��K��z�M�)�[&�TyЊ޲�����3E�ǯS�-�^r'��#"V%UO��,Ι��w���~�|�	g:�4���Q��[�@v%ʹ���nR�(���R���IBO5�����S��j�293aҰ0�Z����N��*L5�7�Ia������?��Y��_����P{���}����d/��7�N��g�>wHa`�N�k֜F��FfIů���kxl�j'{l8\� 94��
I��I_=޽X�(�R��{�c��󣮇�R�1>C<x��h����Z=�̗`mT���,"LL�0��?kp��i4�設�-���|�<�RC��_i<I���.֥�J�U���LeTC����ɝv2��c�H1�t��HI�]�9����԰&#���,q;�,�梳���S,T��V,KY�~ 4�j�!�BW���$V�:�D�Fǩ�8��*Y:��0C�x�;�<��1@�|����y\R�QE+�X܎9�.�42S�1H[M����(G7N�ܐ��!	�����N7��Xʨ��)���{�QIMȅzk�(�Y�Y;0�Ve�8����mn��m��v�o0��2g�|��X"��<c�20Ӯ��G	�f�d�Ge�c=��̤�$ҖQ���V�x9~�HÛ���>t���$�vo$%�"m�o��pAy]�t�K5�J�~��M�[�d� ���h��_���T�ڊ�����o�M��Zs�22
��Yi#����np���sW���=� K��������玠��*<���ta���ަeO��9��~��W�m`��p���� ��4ck *��Ҽ�"0�����,��Wh=C�H4Tک�m�C�O�
����(����Q	p�V(΋�;Z�!��
	�������osk;쌜��̚b�7�]�ǌ:��R�T\�ϋZü��k��<��ΆGS���>L֋�[��d�Y���yJ�Ы�;���%�\�Ǯ�j�/tbl��v`�Ĭ�Z�û�� J���b��,3"���h��ϵ�#��9ւN��^�&l�=V��Cڿq�C~���j�<� �u`,�WC��C��+W�Մ�ێh*�O�xQ~٭�Ѻ�R�O)&�F�f��?=�n���\ÿ��Ż�:�	�+l����FH;�'.jXMH��fA>�_�%��+k!��qXz�G;?a�N(.=���a�*�^E
L�4���Y!�~�����ۤ��0�r	o�z�5�X�N��\��.�������	���P~�(�GIf֎FCLE2��=!Ee21$�����w������-�NFl��3'�+�e0�<�s�x��N���D;Rލ��쉮O�����ˬ�N/2�y+~�W����>q��oCR�����1Ҭ����cX��r��g�t�@)��i0{�Ña��/���:�x���;�����!R{�*�ɖ�٪8a	�0\��:R�("!9n17��C�Y=�~�9m-�r��i�I�K��׭�k�0s�#�uZ����L1�X]�G��#�j빎��b��i��a�nΖ�P��w���@�<�D��=��o�a�K��Swɷ^�tQॠ��$��:��9"J�'�7G�G@�������f�~�(Jx�L��z�-=��0E�����0U��{`Z�e��W�*d���W[����R��ʚ�f�{�����4n1H�{S7��~z�n����f�5�W����xw$)2A����"� ئ��"�:��Ѱ祓-BoL1O��0:ck��g?���
�&
�8�I��0Gt⒲��Ihj���-�"��/{�YR��o߸�����= �Bm߫ܗ����(��c������^�|��%�X��DU?��n�k��
�Q��d"fpG��D��V�c�e�!�j��qx�FP&��KB�˙�厏�w���w�%���=#���p���u��H��m3�$N뚬��?���1UB[-LY�ӱ��)�2k���`���I��m6(��Fu�l���K+wޏ��D$�cX�ID�5����O��ݪ��i�6\&���N��+�}��vfg�Q)]�Jӟ�W�f��0E�5�-�רy��N~�MҌ=*[����{�,&Ԧ��D�|o���V�!U|	9�=��8�~N��tl?�ZM�{ �k� *���z���oES���.���4Q�>��Ht!�.�7.�L��/��Z�[�[�'Vę�B�|�����L&T9`�	Q���^�DF~�{��zc���=c���i4R�Q˹v۟��B�
�ϬșT!g����5�x^���Tx���nyTS��r1�sS�!Z�CK�t�X��<��2%���'/���&�e��5Y�S�NfhZt�=�o�ȩ����MFKJ�1�)�y{?.��*�e=�i�pR? п�h旃^��(�\� ̽��G�p�p��T陯Z3@���]��F6�Z8��Y�Q��I�$��mꂆ�3Ǻ*>�s/ۡ$���7_�5�DO���v?!5$`�H%�/���bB9UK���ʰ�Jx擰�&�"&�$�2�[��:_�ޯ�{�zb�p�,���d�s�~��-8��{�=7�&)��pĿ�-%���I��|�#ؔ5E�גJ��C_���b�̗`-ſ� a���n�XS�Ґ�ϖ%[P�lI3�Ŋ��`�Eb����zw�����P6F����~�����
]����xuV=)�4S�@����H*%���FU-�X�U��8��&}*��nG����m��0��,8��刯6aTx�F��%3ny����Cg/�V�A{"�'(��Fha ��ʹ�	���k;k	����V,N��W ��Z��"�(p��{���.�|rvU��ik�}���84�pL�Jw@&Ƶq�d2���E�B���ŅI����F�/��L	�fl���R�w(Ldtf�.�����{�8`��P�ގ�3(9��o�nZ=����R;����{64������xH�����İ׉�)R�H+M���)��Jʿ�����z�kl��'v��q������Y<(�H����@$���4��9���g|�|5�����ml�I5�ǖN�&���m  ��
�R0��9��O$�m��;U���X�aE�P\�Q���7v٬��QV�e�^��*��-p��"Y�u�BL�E�V)̥��,�����<h��3K�Y���<��3�Ӗi��H���� T����U&���&)���ZH��X.�-��#��`8�-^�ǒ��@�x+a����߻��/ʨ'��O/���P�@.��P��п���>$�X��&���^����i7����_�>��8�7��r�����^��sԳ������ƅ]���p���0�uI��n��a@/���d}�A$��-q@��Ƀ����ۋ6ƺ+���V;�>�_(��aq;c����;v���V
��!���꜉c���6X2r�Rx省Z�0��i'��~[ R���K��c�Q���C�T�����;�P�ll��_���áN�@.j<���c&p�j���7n��	�=�_c1C�=V>Ģ��y���v�}o�<����$KL6�V����TK2&��^k�
��qԖA��n��	�Y�3��� o�m�։�j�Tt�e
j���"ü��̄�}��a�j��|��Ȫ�
K~��(����=8E$JW��B	��<r�<U�ƀ�m5OG�)��?��(ko�d�c�P9��6y��;��@s��H�g����� �U��g�|zw���L�լ����돗��9�%gl�{=o��4*y��֘B�����1g/��œ�t#.�:O��㳹�X�z��cx���S���І�鋛�W�`�ޘw�jԅN�FާOv��),ɬ$����,#�A�� �+�O�-X-Ӫ���6ll�m!�)>����ǔm�E_�Ϣ0�po��M�>גG��eHyJ�x�9�w�j	��L�F����]��K�w���Z'`sη6q�dlh� ;x��tm$Z��-)L�?��I��O��8�Y��<H���SF	p9��C�U~>糜wT�F�o�^�y�%V�ly?�/@Ǹ�A�2Vk���*>O�x�(��<zP��)`�1t�K�����RVﶭh��C�N�L_�9 8��݊��0�X�M+��h�3�>(�72\�e��-�#�Pl�L+��>��K0�Z�a;0�ۜ�6��k�O�:3����.7��^�@��Me�0��2����k�1>Ւ(��BN�nQ�"fկ	�������Q��jŭ9�acF#���P� �=S������}����i�q�Fr"�z�b8�*�Z�o�C?��a!��d�,k@�ɩ#�"�6��ĮF���n�g�� ��`L�E��t�1O��PiZ�M��g���t����ӑ�ﮢ��Ɏ�IeV<3�yՍ�E�'����K�le+r�j�bi�w�D�(�A�� �.�#ș�S�"�u�w�8	��tt�AiO�a�3u6��3�%x��e�B*I�zz�0���kQvI2��vb�h]>$�};."ٍ��	)�
mĬ*����y_9�|���[uTʒ��ΐ��s���W�F.���gkm{	������C+���\3�A)D*��>�T�,Z��hl?��G
�x�w%�N6=y�ZІ���㰚�6�_��oxp��b���0�_7��V"[���(��w_C�����c��l�Ȅ^+L&_:,��/��>��5׉��A�� ��Wx���?�R��]�2�EhDe�m�D��:g�ݼ"�g���óg¹�qK�����;h7�b�1�jyw�Q!>�kq�ѥ�9��m����\��e챬}L��
��bk���})����q���]�	Q�6AL��q���y��I�V�m����_�n 2e����"Ɠh0��^Ԉ�a����v���TJ��4��v��gM�x��YL	ˊ[I�Vtc�,l�qQ��Q��+.q�
�UY����������Bߞz(���	EU���a*�!Y"���6G�$�D����8��G�����
�r܆Ӟ%i2��m�
f���ۿi�X-�--�����O�0"?*�x�^�X_"J�> ��8��!��a�k�ܷb꣨]�1�����+$�i���G$:�n@��2m�r�������Sh�!g��<�l��C�:�i���?�����w�ݻ�@����}u8k�ܫI��E��M�A�)�o��2X���N����:�;+�Ӑ��ՆO��XI�I��p��a '�����r�F��N���f:
�?��D���1�|#~�kG	&b�����������wL}��J��z�&�q�H��.�n���m��	fy
R�Y��	>�4H��[�5����E���ǘ�s�TBuO�+_BA��(	�d�whKIgr`��XZCRT0%���Oǝuɬp�뵌��gy��-YAnm�Z����F��Qi'�^�/VR;7��-xH�U��N���V�VG�o��	�$�i�n�k\�,� {��T����3�VOIT`��O�G������FF��B��!a]���&8V�~�zz���'�Pwo�s��2asm�b6"����/$yVy���A���:��c[�^I�b-�R���:B S����_�<*��#i�90T��Fɑ}/��G>��"����
����8WT�ûJH�c�k��m�(���&�p��ܨ�B�?QŇ� �$g��5�J6 ���u%�x�T@v��w�8�(dF�f(��m�
8e�2���H�]׾�>���X�A���:^0�7R�@��bg��"w��$.��C��!@��kͼTXH;C��$֬Y&��\����~k�j��"��M���f�0<�BgYaBR&A���v׌b9#�%�_ص��+J7>5���F
�G ��/)D=�RdGW����(����H��r膹HLT�}�S��5������)]3���?� "U�+��^X����o�o��o��k"6qp����Yp6!վI�E&���p!-�~Wd�\�1�G3Kɓl�ɚ_r6qG(�T�������J��sZ���.S`�2AN$��;�(�b^Y=OH��:Y���uj���^Tf��*fT'r��.#�i3���P�l��Z��+鋭�#LuI��M�)�>�����:!�_�c�	~�L�8���Z���"��a��(������;��_�e��]��snoE�W�>-W��I�Yht�q��M�ޢ�;k-T�/�a�Q�_�C4�;�+pej�ª����;m"I�LY�F�(!�란y�X��RlM���O�,���Q>�H*ܫ����c���j�Ș�GG] ��Ru l�eSj��~PF�l�c*W�^:�bU@8����<��_h�[.��	�ļ�Lt�ʊՐ�����X�h�p}NC��Ž��*�|����YA����]��7Mjq,��d���BiBs�(�.�G����EE�&���{���͘b3b��Tn��AjZ4Q^�<�XV�OE��/6�s֭x�(����	S�P�WM�*��V}KN��{�(T3d8i�,/�a9#b�Fԟ#�p�B����A�H��I��<\�(��&�zx�$���P��3s��VK�/���q�j�ÝM�xQ�+�>x�hY���cX.�fRLwMBAϕ�-��7K;����nr��W��d�^�rP��:�%ՊNUx�,4��0"	��0�,�]�˳�&���0�Y,�� )"�շ�a������=�XP�����$=�'���l_B�z�O�
$x@�5�mf=��i��
#oݭ�ۛ��4�+�٠��!n�j�VÂ&Z��qsU�Pi��/e�uF�ؽ�3������TR���Am,��-b���;]榭0_���;��\��5���	�s<��u8T~��Bߤ�38HcB�!S)�U4����*���R�gr��lL��ܳ�"��|�K��n*[W��A��WV�����q��N���.j�msr2�?Ĳ�V;��^7� �l�V����ķܚ��v��P�ɇe�%������f�,
w�-OD4,�x_�p���;;��a���4z0GDkvݬY!֧�|�H��咎������g���:x6Y�Vd�S>�?^�/)�5y"�ސ����W�Zv��x�`�@I|~ڈ�t!�(��k���/rkX����U�M�&�ix�� ꙳~1��в�����u �Gj:\DH>?�L�R�s<Ҫg_q��͑Y��2Ra�wn�5I �������%j��+v�M$�~�F�o����6�Wv�����Z����!4T �&���eDe#%W).��E�R��_����G$�k�+@6��
��@rj��'�
'����X�����'{�$ꢣ�\��60�����rQa���C�a�U2%�]j��Q��T˼0��=���U�?�]��^@S��Տ^��׃�hl�n��+`�3�|���5.������bK}.ki�F��E�� �X�r����⾲Se�� �)R|BE��zVH��1m�֝�j�0`�w�Rm�b7)���Ɛ���/�1��x`0E|�;��$�s��>��)����F|*G�|_Ѳ=P�^�]
��"�`����S&ɒo���t�v�="H�h�o��8 �Ks^����(��\�e]����آ�����2;�Gn�����b(v2Ք�ۗkH�2&��A�l�3$gj�V���:���A�R���"��	����>T�cy�^��g-�fT7+B��Br�r��և(U�� ���6��cb�t��B�D�U~�	P�EM�kF�麽���(��+���3j^�-���	��.yDX`�mo.;����oH�JW�K*?=0�:9���g�"bU�׏���ʦ�5�3��H���~ұEG�k�6NG�e�#�H�|'؝"@��zx���$�m�y?�R�SL�z)^����m؆��y͛�Z�Y�ȃ ���{d��8F�r��#X������2�8m�y5t�k&� 񗾧�E&bT[��o#��x3������7�s��W8�;6�(�����̼URu���ܗ���Q�����B̾�%�T�ؖ�ӊ�Ë־��(����h�ґ4	��>I��ţ������4�j�^�_g(�|���!�;(�.B��`m���1�&m�<0�ȧr�fȶ3e�D]Ute��%�F��R���k�n;�g~��r��y�P!��%
]w4��G��ȶ�va��I`� d���wϭ�PA��g[X��Zo9��贳��2�35�K�
��ۨ?3.b�Hk��D<]�6q��
�;��<�7�֭� ���D�\J��$fފ>;��~e�	�y�&�&�-�KWN�!N���%+q�0�5v�_��MԐ��J��	�u�D��c5�M��8�bVzdW���W�9�?����2�lZ<p�'?p�,]�7�p��l���61�*�&�a�+������LH��4ɵ��;�9Q���s�^�:a� �Ⲳe~Wy�g�� Ƥ��@ͦ������r�a��[N͵�AW�e��N�Т��Jt|~�۩�j�a���Y� ���"����%ʻ���X��ʿz�-p�K�)�(.T���M���{*���@*|[�o���U�����
�7���x<�Z�{��F����W��י}��j_p�?�sV�A�VVcc� ��:L�SG��]bP���DF���ݒ�ʉ{�3�Ԛl�Uu����y�ʇ21'ز�7%� �L�����k옠�����i^Jdy�rI�u�_�;�	}�ş���0�:��M�7q3���Y��:,j�8���,�qU,r$3�zbݏ#��f�~��O�{k�s���QXa�\аW 
��g�!�S�W�9��$v�='���k��_.��X�����H丐"����]���S�6��p�"�"��tFG�)��Ӥ�:}aF���;=�&�S>��ۍ�UO��&PC��Y$�5Q��t%kQԯ҅���K�ru�1�U��s�2����J�!z�%s��I1Ϳ��!��P+�l0� �f{g�o�p�P��KI�(k���Q~WG�[\��le=-@o�������{xV�N���k���ld�l|l	i�&Q�ݸ��[� �U�I��j���I�i�7���'�X @����*o&�sX3ɠj�x$Xg��M$�g�f;�ǥb�'�x��%V���
�M�%���Y��{�;ص��aY�"U�a�IAY��S��K;^���q�cd�*o���z��S^�� w�I�,�V��_,��(u�a�P��)Ò
�[�����xX���@:���ٮ~�O���~��4q�E��������vA�r��T��ň{��)��Q�5/L ������s��c/0zj�HZ돍ɒ~t�1��y.�=����1�,R��K�6���?���@��@�B!4�����a8����	u��j�I�0�P<�����t4(�*n�%[g�K�y��ApE�����#>�Fi��֪�,`%�c5���`i�W��k��)U�T]ԲX�O�/ZX�F��2?P5+*A_K�iT����2��wJ��r�s�.���_싏7G�]TȆ��jCw��0������( $`o0j��v���wV%J~��ޝ���I��
����c��?�6��Ǔ��kSS��E&��;"�-�a%ٶQ���}��c"�}�~'?~e`?S�ʎ��~�ΕsO�Nv�h�`����+b�Q�!;�U�PT��k4�IrJj��/_�%��fBR�
9���5��_�ӿ �Y2��[:1`C�N�}�k��7.,�8L{q$�!��ת�{S-"!<~�w��@�j��U~�FP�WW��KY�1{��J-�ӥ�Uv@���ݫw��6�����$u������n̺^:�Nbp�|� �cy�lϱ�yb+P ��CΖ�mC� {��PS�%�؏�S-���I� u�����m^eσ��$j8Ax�3�u���=�(@ps���V�K/!�QL4Ĩ��Ӗ2k�9�Y,bo�MI�;�+|��X1XYN�]5kM�	�Eӄ-�hwW+܋�v=D)<��Y`�y�rGd�#ϐңk�7?;�Gߺ��&Q�#�)����A�q��Cߐ;�-?��+i*\�`G
�r}dw�� �X˘�^��kf>����iRLY,�+7;�r��ǧ��U�$��������'{��c����*�H�63x�R�Oy�#>(M�j&8�'�m�Q��r,�Y�{���*"Kw�)C��pH�r,��N`q��QB]n�ͦ�ZF@�Q�Q������9{n�mZ�7>;1���	L�0L%ս;m��*+}U�"ۆ�
�!Q8�	�a~ߙ��u�kӧ��`�5/ ����Ŋ��5�IlҠ;W�a/�mc�F���RD��	ͼ�u�4e������H) _��Ĳ��BfXck, YI�'����XU�}���V����FS-�&2���B����>����������$L�?ğ��?ˇ�h6ӑ��/��	�����H�,R`}ұ����/m7"H��SЍ�G}��@����|#�o꘠�!5��,�Z�R8�*�a�r�b�v����ڳn���f��"��S��]�w�g��=@���?��E��J���mɮ�o"vO���ţ�VK�[���o��c]p���GcQ&��U�:3>iI����E��J�Eфҵwnēb���9����S$��O/�%�b�")�+ś)�ÞM�	s~Bs�����喋ň����������Z?��0�W��� NY[d>�����$ ��:��!>�P�\�^\��� h�����%�( 9<bM$�>���W7ӓ������zҙ��Bvg�h�#GI���z�+p˗i �>Ø��^Rx=�~L=�^^|�C���^	읱�n�����%���W���	��x6Fim�u�)ws�Z�#�F	����_:�f��.U���|O��D��cA��3r�[1�k�HB��0��Pѱ�A�vx"힥�[`�+*�<֕6�7m���m�(����Sòy+S07��N�q��E���jǊ6�pM���l�r�O��[�l�_����wD[/e����f�UF�x��M����C"���l�e`�e82P@:��F��a�5��@	Cm���Z:6 w���@�\��u� �3�;E��<A����\-@d72��e�Cr�PZ:��_�S!{饘��b!)�g��bh1�,�ɦNG5n�M��sE��o
�|4���K2�~\�Z����HOK�hڍ�}#1�vz��t��"�z��nK�\����-�e��sńŲ8�#��n��d"��0gD�"1O)��|�e��A�����R�I��%'����7���V�9q��'B����J��2�L��g���9��?�`S�Ǘ�Z�2d��'9����X����aRU:��6���2=�
�v�|�Rϑ�핔��@6{|^����?'O���_Pt��5�A�J������s�^�Ƙt�jׯ�D�譫q��bz�Y`���m�#}�����op�":�8qt�Y�ٰ��
':gb��Db���`&�������eD���z��ىdи��PA����7&��̎w*f'�t�1?!"��?��$>��'�;�?j�M֔���[��_�8_�G�b�'��>�Q�s_p���L�k'*x$�̩0[�PsUo@��)�Tݽ]�<1qbTH��=�uDy�X_]�dX:����&���<�n���F���]n jA��&���jK�`��H"��O��]�L��^�s4@'�3/��D�S�����O��p����n�.S��ۡ�&�������a���h�� ��{/���X��6 �%�xQ�&�鄄ҟd��r�hhFv@��QÅJY�?aU��!Q
i�P%�����%n�~�9��z^�?�[����}*0���Հ�G�3�'��ŵ���I���Ɠ���xg�b�|��K#��-�n�M�)�D��i�P:��������[�0 p!ڛ����̈=���(�ĀK̼��R��ݚ�O��W���yL�r)J��̾�T�����q�œ���=�yiˁ/gZU�H����(���'�L�X��������F�r5�#@l��	����m5��Lw�Pl����'	e� ����\���Ri��RXz�[Q�A\A�г�In텸Dk�|��$;6ȴ���Y76O�R��ں�f�X�f(����Ԗ�o��ۭi��[>��߮���"�'�{����܄n��'�R�%?�-Ե-�ʒT�E>h�.���E5v�Mx�2d�nh�"�
,��d��K�o�9U�W3��p���z R�84j�ve���㷕?FR,`�B�Z��sSz�@b�S�R9�ۏG:�AM3��Lݟo܆S!�ɣ ���/�E(�ɨލ�����{@H?nk����\���kn.[�J������!���p�O"؈^u�@�U�7���O�YV�[����w��,Ij��@9Ma�-�N�*���)XKw'�ė���S!�*���rս
�G�(#��c�u�;�w�_�<�?�Ұ���e�.�#m�TG/���2b�_��L��b��@kM��]�T�ΊM��s`���D��c��R�u�Ojs��S~@>��"/rʞ�K.���.��R,�٭�in�����@���ߞ�J$�;�-�۟�)�DU<������%y��f��DnRu3�]q����Ӆq������	GK�KG�z�%��'�$���H>j�B�,xy�jF�R?F�� �2z�T<� E�����!y�5�b3��T?��-��)�7�.�&����"����P���![�%�XX6<J_��c�94 ;�-���m6��h�� �����Dg���,��j`�+
y���%�Ca�	���}���1�*�yŇ��7�P^�P��H�i�B��Aj�_3�K�d\�����x��i<�/Z�,&'�K���J.�����4Ei7�љ�ڪ���e@m�_8ROЪ��ڃܼB4���E4����<��Q�_�M��L��U:"�6Y#f���AAQ�t�~�C�o��J�!J^U������-_�pwb���<C(BM&W���Z���� �r�0J'�������͏~{m�xh��ϛ�/mi)d�~>�0îQ����A��*yy��r��ҋ��Ca���B#����t�t�����]��dF���Wï�m� �T��^����4�P��P�?�-���m��<v�ސO9�4�&:�&|/���������_��E�u9���f�6�}҇F���*�����7�W�������J.���=��@0P�3����zxW>M�!��{�����=r\�����{��u��A�����X���ߍ�<i�@U��g�r�u���
�lL�����^����<J��,ٕ$H�ۓi����K��4��ݼR*ݻ��s�{����N�ѺVt����F:|4\�A!/�E6� �����	2v�qIآ��*����յ&R��\�(�Q���E�6����a��ӂ�xWӻ�Jп�߽E����yjy��̪-�M��K`�	9ҫͽ��� ��v=�K�+�!�j�N[�l!Ӆ��{���]�[��_ټwJ������U�(�@����yd{�@��Pv�ǉ��ղ2�6��i���zc=xE���:D�q���mi�1�HR%�tLmz��P��)m�x/�WV��X�HK�`��&�Eʠy�'$�	��!C{5n��P���D�*Q��@���X*�K[�}:��F|�
j�6ŋl"?g`XŇ<Cb��J������z��{��v��!t�颠_�No�	�~��4���v��.<|=��'�9���U�^�$�LU�Mt�I��\������J!d�ϞίDU���4��OSHO1��f8(b����qE��@������D#�ٮhKdb+W�y�ǅ:Z+��9�*?�_ˊ�������s�©bd���z@�ye'rg6�H��G,L0�K������S��t/��<�"1��i~N�X�����9I�sc璴gU�k�Nز�=/VjF=��b�r1�0N�u���[F^"�wmz��X�X������J(@�*�>b������)�E;q���4�O��t�X0� Dk�c=^j����Q�V$�ibC�bٜ�f�#���t�7B�TC(Y��w��O���D!	Ή[N�����R�z�D�-�&x�� g�_v�p��0�6e*�ニ�_O��u|/�M'���&Y֏�-����l(o��Φne�9����M�Q5���j(��4����o��{܇���`�J4P�F߁�U��c~�5��ĥ��_��.������U*El#!ňɈ�Io{X����� ~.k׺{9�h���nQ�}k�lJ:�L�lɴ��ssαNt���2|I��w�7�(!
�n͓p�g�2U����C�_C 5� �`�n�%s�)f����bO�����gjaxƨֹ�b�3[�7
�j4R��q�9��i�lv k���D���L��@r�x\4�D8&9���p��X5��i�-��K���X��^zw�W:K�)Y��"2��S�e_�P;�"��O�N��sY�?|4Ԕ��.��аC�!������h�*��F79��J3���wC�b�@2PR�y]��I��j�v_�������s8O��˾D)���6q�*�@���C1��duG"t)uG>DdZt)<)��2S� O���y�ΰjk�O�QVOJ:��	=��q���:������ޓv�q���0WfGޓ����w~fgT
��W�|�7nP�Pj�k+ޔ�f��(���P�g���$"� ��ڀ(/-!�c�*�/�O��@�{V���a��a�]qRH��ЊHzKg�j��<]p�$]�hW�d� �)�Z����J�2>�k_�ŏ���ϔn��MaN��:�lk�BCM�s�i�Nu{�J{��a}c-�/d@Y�*�nzR�e��'�>j$w�A����T3�[�zi9\����{��-�_�5��"��L�R����1�����l"mJD"R�G�sV���ٴ�e9�'�\a��,�1D-�H��9#!� ;��Q���x�|�T���}U<4�Ad�)9SD{n�3�ϟ����k�+"\��8j�w�ZQLdhB	  �lw���j0�L�u漟;��~�ݮ���Xtȿ��b6wBY���[H�38�35��#��&�v<��y�W
��U�+˥#�* Dv4X�M�-߿<����]msj�F\���08�:��w�>Yc�K�#��XTS��pT>�tJ��`���C��W�ļ�v)0�}r�x��:���ymmg�2K�c�1/��_�I�(&��Ghf�*���.ei�#6�-#�����k�E=p��R ��}�eh��#�5C�7]a~8~1��̺S�jP�Z���5���/n>R��]�K��ko:vzZ��n�h#%�:�����s�HۤALK�g�W�v(-�NS̈́���+q|�q!4�ִL��G��?k	�he�1ݛ){��|�x������)����Ź�	sm�Nvfcw���`)�s!�oB؜�bv�0昮���%�q��b2��Gk���C� ����j�T�l�5!�~��߫�,"�_�r��ZA�lйb�0&���Qm�=���^��5�zg��A�Q����L�a�:��	q��c$ǜۏ�a&��S���8P�6��^u�[-+�f74���(�j��PL�q3��(2���)�"�}����4��{�H��L��J��ы�[�
xyi{�P�x.ګ��3FE'�Q��;��B�/�֘�<����')��ZM���0G��H��2�3���)c�)<�C��� 5�c�`^g�`�M�w��+Q�戌x��H��a��{@9�G\d$��D�;y�Vf��'��K)�δ��>ZI����O���W]�Y���n-�#�ۂ ���Gü�p+Dq�:���D���`�J���'R&g��*���s���#̞�7H��FV���X�_n�a
�b�3��r����C^,kkj�>��"k�O��01�U���rP���-+��@�5�c\0J��m�.]���t�O���8�ʦ�Q�9|�I�颻 `���%w%Cɉ��q�%�f�IO�c�'�CY�j��f
����Сy@@�Ĩ٥��k^%�=�_jݗ�!��~�"�L"@wOfd�r`=B�~�e��-lc'��φvPYC����2Ǫ����������5L�'�j��b�)�S�I�\�"����H�ɥ��_��|1K4]�U����D��d����n�]u��؏�_��Y8.��Ye��A�|�[N�#Hu�(M�{L"d��e&f�~�ҢP~Wr#,���C�.��R!�������D��ⷼ�y�{}~��W֜��Ϙ��ڼ��g_�:�6�2�Ƨ��{B���H�Q�6B�k#CD,�}dK��]�j_�)c8�����[�"TVΏ�	x���&���a��`�_3�~!����	�jY�d�bP�grW��3�ɈF�M�{3V�i��� ��^��] ��	c~boSs'ٛ+��?ٞ��F��h���y-lV�D�U0�iW%SĿ(v���*H\8��Z��{����J�( ��^jP+.�V��R�2ˇe-�9��J���6Go��mJ����E��n��eR�X"o���(�����oR��g@�� ��[T�S��9?l���0�yk�>�e�:�V�0|��}���:p<����Ԋ��ePx����e�����S�*�왖%��޻���c5L	`�O�e^���g���Ą�"�e��6"p@�����s���rw�����&� �ɟj�H$͒���խ����Ӵr������-��|�̍��\�8[�Dejh�T6��$�����5�-R!-��22��#�(���_xx�+����������'��7za�e2�C�Dy\���0E��b7����!�""�~=�mmJ��m�¶ٍY��`�2]�K�ba���i�48H�cxq$�B��@"�o��l �k��}_B��(]�3Mhf����X&��2(�(���YJ�)�r]�e�)������.�:����6�U`��;5�IA�����,[�;�� �`�ӯH�������ܶl�ƒ�Z\�"-"��������=����V�䶻 ��o ���+v��������i���
�[eF�-������ ��u�q�u�S��k���NJ�=�ޡD
7�0H]wܦ�@:	��R��ҁA,t�;��!�&�'L�(�h;F|��䷖+�^f�P)5��>�WB�QL��,\����T=z)��|D�� �&K�;�؝��O	� -"c��-��^�E׌\�Q����3o#ϭ5���əܬ%���R��c��~��&<��|���[�: !���E�\gA5��}�Ɂ��]�;�u��!��Rҙ5#�q[�`5ߟ�Bqy�cq�������n�wU����=���#b������w�CL�z��hPYXɍ[RThj7���/o/PR���2��~��뽙n� Y%��a�J����l��µ�7%���Ф��0:j����}�P���'�]�R�Y�1��{$���f�%�N{j�\����9�(�Vo̍���7\��^�@�����p?s3��O<��&:фG�IC3�/Lԫ�J�H�?�Ρ��B��ʭa#�U5����h�T���p%��J�P�$�)hI�S���H���r�8�S����t���}�t��*C�7Rh�p���@/gE�ƙ�_x�7�H� 6��J�8�!�R�.�h�UF��ʅEBY(ʁ���'��z�t(�͋ �j8\�۾N]\֦@�����H�������GR���,�;y�l(�L`V��!�B��vL �\��0�_#(j�2j���adJp���fJec5J�*��C��o������GU���M������R_�>��qWe��Q�B�v+%�P��S"��)$�_:^a�,*�P{��)8��FjVH�[6QF\��h�3�I��w��y����4`l�dp���X������%��Zl�G����M	.�Xݚ�OvՉLnk���3���œ�^��8
ޱ���4tV�%��"���8ER��;Ң���Z���1Ь{BK�:�)p��J�z�	k���gPO�X჉�*S�N]��=P�i�Ν)1>��x���Z9�^X��Z����Qf�(�Tlc������q�^����LJ�8�q#\�E�������3�����K�G�Pa��Q�ϼ;��&״O��J�hV�{��0t;�Hk�m����C���[j�k��b�?R!mn'������(��o6>!����~ܰ#��V���!��4�!�������+1�yn[w4��x��.�١X�~��,Gl�vVk���Yu/���	��qµI�A�pv��ݚ�u�π�2N`����Hj䵭��Ԕ���cf�^���$_'Ps�X��{�4�@�I��j���ضh/�_r!�C89q�5G~�^EQyC�TPۉ8�e��	_v���3_F�b#@n�a�u��K���_P�ԫ@�`��I�5FYm\�Qh����Nr�<�w�s^X�z� W�t���'�)ڢѦã`���Ml�O����(��l࣫��
?IDRN�@i<M�=�DBz�8kt��X�!�eDi��J����b�౞6i�$�Z��	�s�ϥl�2;�����z�|]�x�(�K�ٷ�nj '�z�>,c^q�/�+�����~�r�8$��qx 0�k)��ɽ��Q�@��@�0w��r��+�n����g���T�w�4L<��_��|	j�С��^���3���$(cz���)����Cd�p��za�U��3&^���S�]8?��i^@	������漧Í+?c �]�v�չ�],�ɹ^>΃�}ԋ���D����@n�@�Mq����O-��e��5��W0���\�e�7��I�V��v�ao^�������w;5���N<��i�(�q����f�zk� �mkd�$Ԙx	r�e���pO�ډU�X8$�OW]�mJQq@c��D%��\?訵� p�����[1��`$\}e�XcOuNB_q�\A��<�B���m�oT2?}y,-�W�V��9�w�R6�K�]��8����T��f[�\Sj�g����p��`�?z2���QY�X�}����^=lx���6p=�����O��QjB٫�/	:!���2��ӊ\�y3vzfV���t��_̀@{s}K1�~@����N�h�y)k;�3�sF�&n��^	D���� b!�?9���M��a���2|��>B���E��ȶ�~Ai��g,�͜M��!�I^��U���w��4�;k<�a���6�\�#!M�Q�2f}����;a$B��o+�e��dۊg�����]x���q�t�ڑ�����/Yv��l�/} ���YD铄l�5�'Y�FK�+�Md�}߿3��̷��)b>���y�����R����8ڼ�n�.EM��@wP����{�mk(�F��������u��1��"�y�w��?�
�K���/�x�=z�K?Й�Ğ͕"�� ����$��a�D'�c �Q�(�����k�/p��/�?�u�'��\�POZ�½��0�w;6��"¼�M��82�Z���s�ي�v�MJtI�;$���^��