// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
mNyQdnmXOYM3HMFJYD6viu9O3NAEfpEHFCb+aqRGjWjYJ5t3vkyHl4MIzu/JfV964H0xmfPB/0Me
/Y1fKOhAvZ8EP1CBrP2297VHXb22S71v48uqA30V2cnB4LY7IC+pHrh7BTXWeyck3Aw1Y/Oz8PDe
buHr5e7cHQpspGUMvaV0H5jMcGJzBGxTzE1vtyZEeyBASzah94nvBdRBvqn7sh05vanSvJIK0PYw
TzbV8Oiw9fmw4PzuE3F8c99mbEDbwkPO2EEyyqXNdku46wlLkrTX8wbKPrZSTYFHLPIEm4nqqTUd
bhfm5FNW22FEsqiTLNsVb0DF7mfp67RV5Mzc5g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 21056)
5Hr8rC1NVnzmiMjndFLG9szj868738MRA8zU4JQVdKAuTR3lrVsCJnHLZJqaEWq1SgYA8iwXwVb+
nHjfEPqEQU59/32kLyIzF6BzMB5+3yBeB3PculHSjvZOOlbEKvh8nru1K83iacLUYK6RN387DNS2
IM4nm5t3FGtt8+cfBLANPG7NrORO6P8JQL0fgf0A7QZGC+Odt3+VzoIF/wlCruRi66qH/d6ejI2+
fe/XE8dTXOznojOLqJaCVqbcvLWPzEgeboF2VmXw6dYGo3T3Aam8ae1ySM4XTyzwJiW7GIdPnoWP
dL2kd9cIsq8coqCpAdocSLHFBxkwroe8tZd5HM9d67FLvSium0mDjgln0KVwRL4N/uYUUZqsfIk7
2eyY7oBCcGoO8CDGeFNRvRRXz2f7yYWI5j0nH2zZBXkgPXXlgokWbumAhR/Zoy+oQXpvX017bU0h
VqQJ2RoPSFb0nCvqdu3zy6pToY6CtRQxplMobCpHYDZINrAv/H94jQVoOWbzeJCCML16XGnDXObQ
nJWCqbe/2aaTmkUPrubr1k/cxxiAcDUqRMORAcpvgaVnctsnMKbwYI08xzJNKvDUSsHME0sAT2V1
m2uzlZAkVeKRBEikGSRT0YTUqs8+UoUnf3If+lxWqvdM73LZ6d9+nD3QWyaPuYhlfJZ0jNdvoCEq
YykNm0hM+VuXWaNX+B5983D81WXrDfbzFlry/x2PSs92pZLyE6k/mgvb/8Rv6RX45Oto2U82ippV
mQr1+ewwvd5fcpGOL+cOmZbRobm2iSwZ6gpzNeIwuAeiH+qyoeKtta6god0HmXV5Y5V9O2sQt7LI
zQBcwDf11D0PoFDtXNAZkAsjYBWRlwdlp7ZhaqQ6pyVVbNuU87ZQTjMWbgWqBCq+j3A9mEfEvJgE
lYJLKBQe0H1t0lXNK2JR3AV4zsLRbuxb39cW4FOJRF6P6rxt99uvHptmmBabQKTABPpUIbEUyGw9
gx/t41a2Wj0fd5plv5IjlqcphogFCJ2xIII3tD3anWxlG7uF3HNdFGZBfcrZ9kybWX2Xk8whYfcW
F5x2pmfJMjQAgKNqwqATzs39xCP+RvkHBFYNF/WaqJlrzf/LGwr5ul1Gpb0ZHdP34Nuzh4rab4ky
6uZofSxsXCNyAoBi78p7XXU69Zv01s75TKhFUVik1qiv8e+MiyYTVg1wtKYaKBR7NPeoWxatfsHX
mekPMpENwm80vrMTOehFW2XlgKbLkxIBkr4nb3M1Q5ostXZ3+HX7hnGLpuNNeOZBpIJGK3tRf4BO
2rluXJ0EWirpritAWZskeI+yalBsaw6stp3ANTw/rbqldrjy9/1iu3scf4wCTYO3WH+9KliHrYw7
Fyc64wEzkvn/rZdaMmsNoacxmpRVIz9nO7BnA3DU2D87p37SAa5E2p5zS3A5jZn24OGV20PgHu1s
1E8Kk31p2WA9eArYuGaNd4zkA8p8SZLWeovnysADznDDZAG52BpBfZynLsgFE52NyM0TI/56EkaV
5bJyFC4BxCncliwSrytq4kX0Pl8BQwbAwGzYWITqzojpYJ7Tpyq8G4WCyGZhbg6qAnaF6GlKetpf
S1zp4+8YLrPom8zEDNzT+AbYippzi6DvFe4QMcUSksiXUVIonbadZBcg4HVezaQdcpAckXxVUDSv
/qcgFREeYNs+TIqlKenARCwhSVNn44tZJaQvWExu/oQcdY1PvSmR9qM4ZiTPa0OCy0bpt5tgUvIW
TyTq1St9Drh47VKezUhlpt+Td1aW27Acg6NRpkgNYjdYBj8Fb8E6r0uJ1n5n0u+94tNOtdnoPYPA
auHOt7EpeK7QENYuDmcWUSyqpz9cP76aGC2J8nOE5QSf1vmcn9ExWmmuiIzmbB97VhjWWuNVHHEz
QVX5RVlQobtiIJHw9k73JfElfx7oVNXP1K/IlkJDFPrkhqSYd6nI1aj9MiKN+iCRYIDYEiWgqotT
tbCAe6pPPPiZbsl0i5n5LaR52hzcCd1oxe5EY/YfCg28o0T6o9WSmrY8ClZPCs/+Cc/WsdRrSRCW
hIaAMEgqC3jUgWbP6mCk9E+iUJZ3u7mJAaHjnB0cbeuQjx9B+OiqvgT5s9CgaEVRlUoTdTgMpkBB
bA0X1YoXhfbIGkjkDZnD2udMIA6hOant2B5Vn5GqlX44NeUbf17obI10HJ1zwdTaijRr8nuZLx1k
myY0T7AILwLc8u/FfllsRHgd6UuSryuTc5TnUar8/36ENL0kOFQPB9xvIOfQfXXgaXPCfnKfqqUA
HU1TMz/7dnJiTNHgbmkLmCV6t4g/M5Gi+xvU3vGskzKeiQCzIxKPeBjHX+7Ttkp6lLSuBL4T9THd
pKZnOAq7s9lpbNQbJlKiFkdRsFH9T3Y4q4U7PH+BQChL+ybeB/HhiPR1v8/TyCocH48pvnxKeEvP
zFQNpTReazSJu8yYhoJ9lD+9t5bat5b6egOOxoxMY/7w1Ka1RUmMZWIqYcofMr4V3fqHXooTmeX7
Wn+E4tJIBuPypWKqLSUdJm3gC/XQWj5wlsnl8LDv4Mi/nJJg7O4OSeeNTDcn+phaQTJiqRaCSNZI
6DIjShT32b/bxjn57U+K4GmiYM9DmdjLT+v+SThG9xJrBmh4ngHe9tHyA0midoiJsuBHzPR6mnYr
6qkKzNzOAQV2reVqZs0Gl3KZZtww5op9idDmbg3dWs2rZdLTnW1x3Y9kwQi3c4TDrP54mxnDNLiE
NP8TD+fxmzHNUpcmC6svQv7CJMlc35LXpa2/AUijamO0nWYVWfunrLbTPIBVT6oQoZ5mTfbJnkLa
yyXYWFLQFWH6nlJBw0q+RWU+lLdfzydKcH3oP6+4PcyI2Dk+jR3w4BOaBvOZMsyZtx53yfJLzpDp
cDLcBk0xw5k/gLyfijyR07wrISYfMRDWJ9qt+Zohypev74Uo+uSo/M959xwpJyPL7Kqiq8ui3iY0
hphymUIs7GOLgu2KrNGE+iTwZaKersSLquLh23FUnCtQJcEAbsyAUbDSdebtf87umFuqqKroAwb5
bd9ptLpyvjtTwyhoO/CEb1YUOrYB+wxNUZWcCLF4rJ6ME7NHKtNcdG6nhITRrrkWrxaVP3mlKWu0
VahOpfgg5PV5+2ECEwdZ3znCF3QJ+XoqQjzyWvg+O+8J2Y8m9qf357KxxZUqetRjj4SLU4ii0kWS
HX+ahu5FXxP5zBCfdcIa8v+11Ggw3d9BdabBqwFOz8+am9NU4cYZLHyaoSMfOeMtxqWWRSBTG0xa
R4+7mguYgVhL5OM2yZ0WktPLl5ulwpWL5UiwYs1fKKho9TYQjSFe0iQk2TzLC8QUiHmeEAuKzOjz
mBWoXYIS3oSgdGR5FYw0AVKgTsvF85UOH9pkjW+igogFRuMIi6cvnVyXCmZh3cl9RxXUoO4DHW2g
nFOEsVZGiQSEe25i4QlSlf8cZEKXIMhXXZB42+kw1kt5I3j+VCg+lpDx0JZsfSpXpFmOJVmRmuX0
tlPa2Y4OkqqENuZgIzRLsTR80D0s3FRmO9EGydXJqzlWkYaU+8D02oeiQyMCvCS6wTB9ZCmKRmaD
8grlhzv+/M4lqE+OEaVDeHEyWniOu8U6WTOsl9oNocbiOa1IfzMiK5qEWefDzzPtGvMlcDZjhUgP
EzmevOVqjvbC0KrzgZFapxcf1BxBQKuM32jVs9WRrjgqV7IQlh9WT2WJWr5VAU8lmZslV5PqdUV6
n0yfGBRLnLdcZsqhtz3DsignHSvTqGIRHpmbM9xC1Yhg7ONMZtvn+Q2mH8Hkr9tDRzYhYU2wXbJV
qyv92ilGYRn78GkxocgFB6xRV004YewpA33nsGjQJWXcclsMAi6AV8sxak38fTXfdNkIsYlYr0Gy
Y7yDQ0qu8NoIuOWOP7ZPRHJLFA/WPYHBgoqsdYKorlVHT1lpSSvP8wMW1P+X7MD3QP+ToymInezu
1wxJ1cw6/ute4W7koQxilns8H2A5IWGewNx1WCPM2DaFvjrZliQFQqozl0Rqn4oHVf4q1ZerEK4A
7yks4vioOA1v8aMyRqJzyzyf07BtX78IVOGxU6bFrHnA1bNlvxI8TAEDThZz0Y5OC9tRpLIfrrXJ
eQnVlIEQwUiBHEedws4qvy30MX1EiQNX3VRZQqdX1TydbANeTzRyd9suFMq8Mm7XWz0Aws3yTYUF
dm9+kaFE/6NcaHBpBSFrvU8dqirjGtqPJm1YzyOwg6Wb/HDYdazdT35EiSL9p9rA3cs+++miQ433
aknHEb/PcQ11EgVUqk3f559ofbAogeUgna6pXUnqsH39X4p69oVQe/WMjpVa0y93UE5Dd8nFX1PE
neNZmxEMnCTe5/XtuPJKkqbh0JlysjKraWedOZvGdATxy/2k+oMdT+IiOhh2PX1/1UmVxIpFJPXR
0qN5o0CkT6sWV61myoKVNvp0Cq5l/HWFR5a69zH0Sp/gAopcCFDSIU54J4eB/fz4+fGMAEu5kjcq
Lpym9lijhcq8mW3bb0RjR6u+yDBLNsFZ5EkzTMGrki9L+6Fw+ApDjfSj3RavauJacmAqUDOZN/fO
sjk+egxLRd54/ZNwnxptrKvMTWcAL++4/mQGOWzuoPIvdX6S6UbRJmFlKgGt3DWS90iATE2lHWzu
Ajpjd15VIZb1GXkS/f+xbah27RXb/n1g3iOyUaF8hyz5IJ4WiSXino+IZykpnqSps428WNMyqKEJ
plx7NiARx/vEv6cvK9CktSKQ4BGs12BHcOVocgiMbnit7XtTEZGnpXUBABKeiwJpRv5wPLFUy72/
pnjaHivX0sGFI1uX3c/hQuXJz7JF03+fq1+F1JKeAIZvQJZkn+GQiUFUQoD7wQJXczeifh1CEPI/
0lp4E65rCS6d9Er/StJaLi743eFy0ZPQEvHrIPdwJZYidjeWYSadMy9GlwMaJC5nnaf2l95v9jGl
WACOFZtumfStDLwC1O/SvjLfaW0TMBrrOMMTf/nGNyF/9prEYugqQTXTnuKBv5ZpEeyZEOb+Flmv
M0lG/bFyHfdgb565YzR59EopRyCf0c1g7Hse8ZiNbeaeh37Ni3pg+vM7Mkq9rqc0RaZLeChBewxH
V2pgIVuzPifGuJnK2VwwtbK4HaodbVBUNXDQ5BgzX6fjP4OCtZ6Uvro0CiDKlrWUbyeVbE/dYN8f
t80eh/Q3QG+grRcXkMmEeRTwWdtjcZ8VY9amsxtsan0ThxVHKE0FrohPBtJ8fQjlvRRWwrW/TgsG
RPMs64MerivpW1NGt5QiS4lbUexkgY4anlQzqXfwA8jdYhPiSw5rT6fZDoK/Jzd7Gka1jtzBukP2
D0CnzI/5f8RYp8DJxqP0syl8iw6YLp3Ky5aBJjM8JCtx11c80L6xaOLLiDkOady9ibbcpcgnaAGM
gWvKaYM/U3+2Q5Shn5c2xeQt8H/ob0pWv368EiQiF/5p57l2q7vpDnTK59XMRmsYFmq8vNz3ex87
YhQcvzpV7Q2CDHUcnT3Pl5uDRPrnRui4nJKTQGiGc+JOnY2DlvoOsy3VIPFbd31K1LPjJ4uAA968
yg45CqSR7ERzOYQvGWq/jiZxGkt+4hC/ZOE8Wn5aAzRcZ2jULeuHhE1shr7KQrrYGQyFxqltZFMF
ZOXAfzX+2+j3nC+1c5U8BTHeB6rrUrL666Vgp0e8PdsGbHfIlEaGoSjuUUIU4hMf6IBExr5aeP75
/7qNB336YtY8W6WP/2goUo3OmA2p6dvCtFTePw2/qe8CjuESMtwQHwppBEB2sLQT5ME6q92vYcBe
JnQIYKwAnQXWL/ApuH43W7bjevSgY+IW3KNUqjCxP2OBk0biaec3KX/yF8rzDFHuetat0pNrnrHJ
a6bZR57z+WbcQnKdUib+bRK72zch5hPq5oF+BAVUMms+fO6LeFucpQUOJQY+oUy70CoyG8mF8auD
QqFKpdns2tkuHgE2xc/kVtrtJTiIxg+gQ1RTo9mAyHInycd13pZIxBLN6HrbRMos+24+eBAUIf2m
nK0Y1loMFRb/8NT6aACCY2ylvqs5OmQRKO9EGh+ASBhZDkqwvin/WjqhZVNff6Tvo0os+OvUjfqB
bCIpNQvScGYJkwyhCQDx+7h2UquZ0TeSBR4zlMHR+ldqLZHqjufqYTzrifEBWKsuMAhhCbC6SNYW
6T/111sqFHGQQ+HQ49CEiZacCH7QjCzLoPE277epXVM+H+AKYS9qzoGx0sa2vj2s8HUhMq80lvSg
8D7bKxPi5AY80VwE0PZrOsCe3v+skr2qGg65PB01mY3v+OJGlp1+z828dfXcgaYkQpFAaukvLtZ7
JDWWmvQOZYqTQ68lIT/hQhpEV9ahz3hXCs0AYGaMM+F7pVNISOoibN4gIDfQgUGCJ78hWLzNOA01
LDceVa3/7zO3pjMD4sNWjWtxAJRqdQImSsOd/pH28P0gJpnk7MXsYDG5qbAiciY0M0D6Qqg4ZLCh
Iw/4w1Yd8CmP3BHsWQmvUYvgCc09VnWC3llgxJvxXoXlUOUCqLrVnhfQXjA7soRvMNV5XAAFipuD
dVAW+bw1jooxXbMnzs/UaFRnOPYai08XbHqCT78D/S3NOQtkqNes/CQfAGuGKnYtRr/hhvpeup3P
Xxf4qgB/0XSpCMNaPUtDHgVgCIcdJBqGgiNZy+YMwVixEiLiyUM/msYY6C94goYfNt8bWzB7atx5
BXbytouZGxi8Yj+7xuMUVsHqqrF53iIaxdXTtQQF664mek7PqseuKxjufYzpTO2eF8SQjf5VHheM
0xB9uCGjHu9ypasv4jKmHNw3n0J377hunwzSp+K+MZPc8SZszr1iS83L2if0tPvzFDXvif4Tc7ey
V4b8goTZBqUOn7zxzGQ2VecRD8JPxeFsddy+0R1JmG9mcX6U5z9nVRSwtUVqysMt0p4hqJ0MlLEM
VpKcNRa0LYcqy/AGs3zeMJVJD025ZeP+YrpVaUhH6lzrcK87y9zpib4JL8mfU5nLgjzHNSkIKEBd
jZQQPU6cAI2GOb4seiqTq/AGsPmhNH+ZV6Nsa8L4zaU9oouTgtEutab1IVjiSb7OYrFbNw841Tj7
o3VA7oIOyqCJKQdosw7pdfIaOAzt5LjMDteVwAClZ/zd4WpllfxOSC38CzWTD1Ro/bZ9KTp/UyLH
iK3ElEV92lLJP47iNKXeR6p8YrLRMryOc9hbaWzU3mjsH/lDyXU7OxtbTZMRX3z3gAeAJO/uPuiU
Vmfa3nl6L2Po5wKeHudXZDijw91iDyKgXufqgqvGkDamSjyFimgxOKALx5KHI24cvI1r2wMFNM9n
4TJG/bHCRjJloknLFbVv3BNiIHtbiNjcwPWWtTIvvSiP4NrPrLZ/qbSOJd1GAoxdzio5YMLx/Gh2
NzdSV5mT45jNFuU0i82FIBZqkTUicH6sBYFWtUkPS+LE9xytHHrwc3aOKFbpUjqCdNzhAwCoOJvA
mevcsUA61YaGeqAeUv9bbFEfYSVwgjn2kyBTIgvb+F+8f230vPCj9/PRF7+2NDXoaQb/YWDwVsrz
mR9NTlegF9t6Cgqj1EYsgVlsD/T1AAdDTvwxFqMdo7f/ztYBRT+1+zxRSZJ3KNhFUFzwPbrr9g8b
xi/toD7Fgsse7qM+qifV16WrgwFfcB2d5XzNp2fKj2mvJRcj75QT9x99I8ZJkPvoexrGAZTmbWIp
5WqzMMqNBhXDfqC2RcsE03ktLlAOY7m++rRrkePvarRoavWRXbl/oVT8SAq42b6EPAdDuD8CQMDi
15RhWIfaavOzZgcoJFV5y0U8ABcWIPcwK8dGUujlkRceELhOsbtukn6yV5ZifuN1n1pf2FtpZumW
7KzsAqjQxcclv8mKi9yR9eZdz2R9denpv7mG1lbye8znljIs9xuCwuWgyF0BXkoMEHVS/o61dlx0
cZT67gacA8JZmBOVba7Kl6anzgnDajXqMNVaSceO/thwENFC4jEdUK9OXrt305riO2hNKweSVSoN
O8KZnJAPOlOnhI2/NN7+4tVnmUX99aXUs64lLvlu2m1zmCNc6tvvxJ+ICUgZaa+qCFKRUcE/uyu7
r7C+ZIQZ+K4ERhBpnUqyLGDfo34N2CZVULgIWEfhJol7Yt8MqsqVdoFIQdcBmpBEN6pbPuvv7oYC
zCHNyng7GJXbo5gKQobxqed96oPEZhzQz/Ea6z0uz53hpZrObeEsrOibaLB1eQ9WgFfR0qIWo1Jv
MZzW90znddcyrxlvgiwUyVjx8uWElxKBfBURPWHXhFu7TpwTbpwLPl9rVAaL1eAuoOi5+Tha3+is
60Lhz2F66dSnKjeO+GNZom11q63eMG+HUcIxNwfnZaaCNGmYlgprr34S32sRsIx0AfVIMXxAcEsi
+rkEzZ4Ru+/C4J1FJDfE7jAcj0rMgAmG2RUpePcycdJIwzTqQdVyseyGwzYooZo4CykfhgiKephe
74aAx72pNZRquwd6RTJpk0JLlZen940CKoXBqrrxwYbpf3fyYg8DnXgy1oRoxRO49/hKr9cL8OwF
c3MeXJPSKNOJLZut4YTFomVc4u2vNCusR5kPSg0PQkAriT2KtK3gJBpgDlZg3U5fYSrCHHgnXUGG
56oTbLqEaDYc5BbHQDy7fM3+/zinNDHZjYSSeCdOzY9X4Zmf5bu5JjpXzy9JXbaIXvzoTQxuPtOj
CAegZPM9kYdyGfBWiHn32qOaZ4kw3SsBwaZKfl+QWQ73UmKoRVBi1bHfyTP+eJyApkth0z5Qo0yh
0oLtvUQgFFh1x9048+6IIyklk+taBkTXK+7l9ZMkqAaPvgED03X/xRlmEsuVhMLxNV9ALtylhow4
6y2vnZmoQFrIKfQEST/BeJwNd/D5lk8TsI8/MUIMRrEaec1JjWD88UYJAHmAHyhTz5AUnHqdRfez
TnHeCO5SyeIxOMJjNG0+EG7nYfCJhCGaBLaxQRmxPZx7PZ7iMQobc6Pg0elh4r6oMpc4+RiZWtk1
Dxth0fddNPgYY+jxEReEAsrXMt2ZgwaB0W0JoQ7Zh0cZFJrfhRBujBqOCIHXJv0uvhfvGDWaHdwe
vBNYinscJiHMWLi1X0W6b9uJy9pgwfQ4G/CXgqjRdizjEZN7HS2JZ0c/vIzQAOyiqFVa4sw9xZlf
PhljmmfeT6EaKHYy6TMBaN3CyntjR9cb4Qcm1oQuG1wRWbWFCCvhSDLSygYg30JEpaH+LjWm9jj8
XsBgV5C3kPv6eTB+xc0yzG3BZZDUmXAlIyVUHfq1q1m3HC4TLPB8nDkil9g0YcV8JCOX+rXRrXTL
POAuetW0NI8EW61wik89pinnoU+iCDjT+AlLjcSlZcFr6Kir9GjkCCWY35p19iuLaPqnfp1AL/nx
9iz573KSFj1NECGLKepZRe25tPzbOnGDWxC7J8gbLLQepEnNugaMk3oEHl9b/tbmGhviTHy8bMYX
AcVmrj/yuUuIVn/rhtP1jjqYdg4+1Sy/cJm3Y8t4VQ9gDEeP2bkrnp1+mlJhpLYEa7xMQVgRMJgq
h4qxBQXhDjyqkYXNS6lOcdwBcwhtqPA/9aJsjQvRoQxbVicxg3pBggkbpOT+NB08RrOugDHp9k4V
+izCsMnlGNq1QqI1tTQ7e1TPo9wYIIs0GEoN5hvbktAC/8WzyVJ4G2OCqNGvCN6J+75m15y2Khln
bSvps+NA/J3oSM3baVWjUtdoFCejBn3pIKuzd5dRHzwUdBDjOSoxUwbb7QFXxLObDQ76kvvHo8Qb
8QZvSl7eVqaA/BjyY90589Su4ux4JyrWH6nP2Me6dPR2bZsJhP0D58ohAug1958n6qTwXTXkPJuM
7cp5vWh7v2cJzrSaM5SNlW02CdYgXknQ2c4UyylxIYhLTa6SR39lMRwLytb9tdQ1pDfxGsCMEcHZ
heHDMaML4YJkOLK/5MqkppKskkVNW15aPyA5GHJlOYULt8SfSoqAVe4m/tgsMHmEljO9lbfHgWoD
HLjCmjHtGTRzLgXj8C+MuTJ66a2t0vpIT14RlgsezKtPbRhz6BPgjCskTHaU6Ee038TNxVMJH0cI
I8gc4oEAZj0y9imoTsXNFUHk2eEBBo91DKvR0Bd0EEK3GWiljh+zN/TN2YsxrY+3ATXPmtpYT9wz
2Nh+oxEfeSraPCzvcJhejMflVihq53n8AyTWGf73qzCtagS7PzMQCBBnnGb4qy4z3jJZiQr/WAIh
cxckJFgJA1HFG1lh5S+Za875/jK24N4VIRrsw/MtqzXyETHEZoRNhhlgVf7ND5LEVWd02SLkWAVp
bl0Jfodr7YBp6tEsVPvGWPTG795nJEeJNNOJsCUBl2U9xnWqKTbHc7nmje+wFTEgfLvblC2f3BGO
10zbXrZLsKlnzLu8OnD3Y3ttUtywPwEZ8gZaBLqqZkyPAr8jeK62hcERRxXJ3WDQwZbGGH9v62He
XfrmThLGl8KQekdk0ExSIVmMAMCgkDX0Rf8KSwVBPIqRtxsFTGC2I9xmtmmJZ19RCZsMZImScc+l
JV3mNyPbermpeL0K8bukOi8KtwTh+/b7QroV/0Tey9dJ8FmUvnwQ77IJfXmvkOOVp6s3hSB5aYsD
9SmF2OJlZgm8xSgkLHUU1zfCtcdbtmUIJZzbSDARhUgZFaIajx29nu8aKfFJ4rDqXIW+l76ygZT+
YvTtoXulzhK6eNXJ6uSx00XKMp4Ltm2vavw67s/1uVmXJ7hdfCjaFwG3g1tf8OZ2m3SoxY3DOChP
Mwn3FphmQs3A/dI2TPp6PjYnq73EzKWm61aOZJK6Ic9SsrlgdZ5NzscN48yEm5RHq4DTO8W1ZB1g
xWkUui9Rsx9Cdd3mZJe68I2cvTPvuUchuEGBtMYnTVq9VYSxug8A98p8PpRZlY0de3Ewu0X7ZUSJ
HINfdLFcUdth/QSnaqEA/9cawviJtMjFkYnlZtfjE80iqmzUIiXAYQ8zb5u0mRNE2MR/zMB9RRHO
J7r/P2cpbEf9dj37B7EEuTXh0k9JoW+EK3EAp8FTaKXkF+uZUeV4MevySvwMEiy2kmCE1bsfix+C
uq4v0B6UWKPsj3W/1Z4o97myMZRm3qfKJtaFXySWZuHNnBmHcg9RCtbswn55B7yOfYezwqWVejh0
+EO7lm/zghEht25ALFS3dEBxXXQab1xqtUAV6epZ37PsgAl/20gdWyxtI6Ovv/0MN8beISYmQVcM
YY7MvZoMrvKgEw7R6OenGwUFksBFLc91EcVutjjgheOKva6VInN5a5qrgwBLHsgU1fbprUxEQ3W/
vRgxrMH481chQftV8mqWGFY4MhPPcu26xkhYDQxBqhwwx1jYIU7sGE3rfe9a+mayEeOjYroRA/2f
n8zLFy7TmWZVqT4ECfnqxYO/AAG/Qrd2s7DIxbkhg6XlH/A4VwzMkdRbyiNeln31ezErsr+/r3mX
au7/ciGSco/OZ+EMdqbsKOJOiAUkfmxJZB0qSoLNLluI+ma4EtwFm0zUu6J0xWASUlTHHbUXJenK
qYML/NsIiuQv9nlEEVYFWZCtQQ6xrNMimniHvDltrCd9HJAzk1Y3f+kLdEBtjxTZdiNRdIfUWJXF
GiiJqfJcDk2oSuBNzDnV9V/BP3kBWz0YJiy+72+cBg22ZLNga6JsAgVCLQI0eBsd78vGci0odnna
UbKm/cCOJkuSn9gKwZyxnE7pqWvGUCWdPrGh8mSJa6fLlhCjkJDBZL+Ln+SHIsDbEkGXcdWVvUtr
WKKEbitCQ3K/+hx39kATfv+F/0tjCfR5Q7k13zsMaG+H+gGRHuf3f7eNqQ5T7ySvgu62MZQvlAte
49WBGz6S2Yx9oSe98MvQATHcfBQTmTUAeeMCZul7FFZxd0daV3XuwVHaW5ob9TxkdU3SM7pWLYFB
i+sfXtj424olYs1bJ9Zybp1XXS2dYQ0uYrnww6R8XguwmwBy/2KnzE6v6O0sQnABLF3xM52Qkb+0
yNcLR2ZjrCRcxd1kVIh0fNEeQX0stll3AkHdWcSwHubDKGOB+qSeaqpBPxwit1GbvA8vIx8ufFdw
oq++VlzWMtVt1Cx4s89NpiTIv1pb4Cyv9vF+QiPAfixlyNV30xTztPaajeA65vQrLRRPdGnLBAXV
ETiKOz8mvNFCtfoPpHAF9l9iQmIFFPl2vm6gf8R9Mc0AJgOvHyaVs26QvOxYUY0wg10REtAnIX6w
UDpPkO7P/qN+g0zAbUEHSUNK1ioCYt+PJkJuh//ae/uoojo7iaLx0f8SBQXkLAPn5bqAGLUPftVc
JVjMvAhgYdgyWlUjGzyYHkdSCKS4nOjFGAC70oaIOseZQUec/IdavYAis9xj05ryYwovJT8531Q1
pm/Dtpn+Azf/kSLzbn403EuvrhjBCBxWKDSdCldrr3a6Bst0+hd5mhJzweJhIb9fa9NhQpmIcpf8
42oW3iwNRnLMAJmACdjaJeqFDhyJjgu+Z0PBqIg5IQABNR6HzTNnMDa/LTQPCEmeKamq0xHADGWk
5JvfXRPOEx5IEUPsA8kNGCClakvtRaa7qeer+MFsCFrscUQuH1oe98/wF8Shimb6biLqCc7ShSHe
1rbMfQGkVfzP2SXMvBHJukS1gXMrE7B5CFUDFhrG8I+jvhZ8GhlAb6MVbJSJxTBBCogqqIiVbWc1
psj3RRcb6D1Gy6BRplCsQLwZgu5QwJ9ljPDi+xX9HTTjMSvdHPKPNsl32F1ecyo8MmWs7mEREdy2
Glb6nLnQLylRvEkvfhFhUHyYMQIJ5y30O9N1Fr2pTPDDZi5Q+WQRR7ftGh4FZUJmfG0i46eg9iAz
LGeZnPuHr8tl5mlTtRuKVHcpZ3RblE8ovBsu9VsDYZrvs/qAYqTstA0hiwF6kxJvr0znNlMYrEQT
KQnl4xwP62OQdbi5zyPW6kAH7IT+CaM5xkcuMUljAmWm7O3Kei/lsARp35l9m2qga8aDg21jkrX+
bY7axhaPVX1KDbJA3lf9KutkRCyihmvydIJIeeubXiN7Csar95w8A6RWoGXAeROrYra8LokR7dSA
egb5gE4biCD8c/3qM4Vzb+7mawmAnvX4H8sZ5QvImlI5tksBcrxWtDZl6VTyiSbXYqlI/T7y07eU
v9O+u6sWvTc1sW512ZujASRCS43xy2QfC0AAbfh5fHhP8XhEJVgEt1CfXDMv5huKQRE0xqu5QiVL
5aUzWMD6SV2IMsStyqKbYBPPfBAp7+U+Kegu4Lkzkm6vo3NYSnj+VLxC1X4KZJJLUfQEgPLshqV/
TsyBOzWidV6L51tLDz0y4S/3Ecu/Xmo8AX9WSSIiL37nxHot47DAbZOFN/zWOUMTjwyXLon4vOHX
ZCAgxkRgCDuf2CX9w7JIkFMTjXDP3eOtdkY+QktsJ3xqHxt+rC8s7D+ces7mvgzm5jI1hS0rgPJ6
BojF2t+JRva0ZuQPmNren3LzqhHbYvG6omE4eLtJLXkXitifpwXk8/mjNj8RhjUQoaFPSkV3Lp9A
oZth//bWXVBmmPeH7d/suPK+Y4H5FARh6wD2aL4DfkxrbpVW+mcM3PRiVlLujWeJlITXgy2oFgG8
/LnDvP93YUFHO/p99/h0c/3BENBzBkek/+g6lZgxnjW2godk461OUkpv8t1oUIYhtLxHNxQSMQP2
ByVKF8gbztOlBU6MBNqPd/05c/QUn2UtAZL3r9rE1Fo7VYau8FQR6Ex8L06XobhAeW/qj0b9cS2D
EUsf7YPzdDiaF+0sg4J18XtPX/h6bEIrWCtU5VEKPICyCQNJVvL4zzz9E3EpH9xO6/1L2IcccLsW
BkB7N0BzRGLb+ADT1Qlg/P/sxlSJgrFMyolKx7BgLuo8O7mYxf3yaEv7oVAxdVjfJyKL+I/tJH+1
7zmHwTZkizHl83guEWXf2XcOds7TwYkpjZ/SQL11PnFghb1WgKdU9vaTeBh1JdHfShnTUzMXVuvu
XeRyXZyvPoKzh0SpJMA/Qo9pkJwP5QWEVzCO4x02IKiZAb9P6eiDfsBd15m8MaYOdsg+HEBHzGFs
TvhCr/rj0/EOFVZg/zcjm4dQSBq7vDmLW7fUUrnKtU/WD293kPh1fj+uPoGlRC/sfDJClQE5Xnuz
Ecviq/H82DucecSQie0Z4LFcGZ2untwVXhi0bde4QOqFLKB0AjTUTH9vJryzlCP09Dau3xV5GjHv
/nTDCKXYWiKfr+Ml1Op4a75DMt1VkzcLh4qHLv3IeGCba4WhcYIY6OBQKiK8IMp0YTlW57NXlG9Q
w8SuxHhZ2ahWf/mRGCjYltktrUVWywldfDlyPfmMDiYHbWBqb0oKkkotTF5jd8zwXeqGayZM5sBm
fOencGr/El/dUEKJoRzO0K0bFB56rATWL+q/RIy3ckgNLWeeX40HEr9wfnX+YcPvaWO9+XFCMQCo
UCzYYvbYZP9sIQGdM1DHBs9wGt0hNzpOlYeXggIzeUZiNq8or0rJmQjN9cq81oXppd8G91t3cv59
TbKFISY0gfu6w8XdjN6a059ZNihWqv4QG8gVhSv4qFgV3lI5P1/iWKBM0slJDrl6kVwWxeOJMeuq
CSUUBhBh6VIyMg+o7ONGqmkwHydTdPySd9O1ukZ2TmnnRvp+WwbDKC8ImaA0sNmIoRqVeUQ6UMWc
kR1hEnZ+CEh9A3458fJy9+6aI/lRMK21gXSE5v1WZzjNx4iD+H6cYtVudrV2DZOyThZTO+aIJB0o
KrSoq+LY7zSkzRDxv5OHzwrQJjD2XTYHcaGLe8HPUaVA0eIyWb71GlNnq2UFEAuTa1ULnLUZu1SF
ntAXJrTeg0JzYkAS0QAyRYi3PXKVDPBYQ/3gn/kRujep5bG5ZOjGuQs5CIX6K3L5LP8sMn+tcpAW
c9Mf2CfMXUnKeJK7LsIQ4a7RWwCcIn23rEggwysam5uBdXT5n5c50PYJrvkYNe5JmgCrW2VuOGe/
/WaW0I66S3KSaudLLiNQTsQCwdxoNaWJX82kDjpnCqKMX/s/06synjuP5m9r9r/3vORdx5MGirQz
X5cRJjsnLk0HEloIfSLOxk7mwjSn6iIo3nKttg6necoJ/JoPhSURAimxCcJgnUIxWOOzcZ7WdFVw
oEpHtCcgV6avHgUV/Yn0hZbmaajGk4Dyb8dVN4yNurNdCl+NXvyo0grqQWVVOsKLjwYORYpzcVGg
xmZpDNh3hQl0bvvsFnVpPIZMeVn3hgK9onlrHJmJ6nhMyByNmIb/COEMuSPSHVTaAMZGSQuweOhe
Q3VFkLwfLYGwWKNZ7HzH82RW6a6w730IjQ0N0K6sO4VOCkX0uqDMhV1cM3+qN9BPBfqXtcTUu6kJ
AY1QmthSs/Z70lrLpgek/RmyOr2DFrKi1rp2ImKuCTSEpqnHXI7DIaHSpX19ouLHxKAwJh3LTnkh
mmC5mQK61e0tdHaDA3+AiE9j/SE/Fu7rEuUvnOnMvht1u+PRRZSWC7rd/XT0FZ8fPNzU2tTuJcXw
kTvD1Fg4L3t+efILmiMx0/L0qFSy73WXiPoMKf9PJuvqKANL+dSLbDx7W+VaGDVw0QRRHQoFHrie
AUXUn+ZsbkZ0R1JEqqXZykeubyhNcxLtkQEDbFHVKo+pBc3OTToqc2sdy3P7yMVFDLRmoYKjspTV
aP9D8ILLLiZ9/KjledppnlL/R5zwpuEfjOSTxqN+vfER5fecwOeRNL1lWUU5xDRmZm2ooWFOdEjl
CzY8hOCsyRW24vOaAuxMF0uygRLpE8XFRih8BOQhwKIL6sDVyuZuS5D0Zr3B+Q/i1UUeZvhR77dn
rcq/XKaFH/PorgwCs/aUAxQIBC+BHUdZ4utw5m1DHzszMra6Sa1busSDx52vec778A7s71fAAInc
t6pUfIBNBHqg4+TmL55FzfQYNiyYqwlBIS4REzVEpVJPA2qxbNnVntrDB2atNJpblf3gP5FhNk1P
HHHdXOg2Qm1h0szXKGj9rOVbkqiC9eeoY8kfuVZnZ9h6DtTGnmpZofce5VwRQoKbSHjmAKMdYY6S
mM76uRxVyuWJ0segXdTRoAZ8Kjm4SSMBzFEg8f/Ux3/LgeyYcKJuvrq25s36Lvup9nYY0xPaf5kn
hP1dDW4Yosl7cfRa9FQVYQgvzeh7ZVY51+ZdhSY0NVB/Ge5JWjMWT9kyiV7RH2YpHNMvzCik/8MW
V2RsrbFsbju67SMxnp0WEUhIW316okXRpPeHHDN1k+xVMieAiylS8XeuHm5KE7za0uEqQy7FSMDh
lk8MN6LM6t/skmx3UOEGiXySUd3lPFBiwhkByH+GxaBhXX/c6DlBn2e8uf0zkwyRKEax8vE4ALi7
8NMSkXw8Bf92RcsZ/6COzfUO1Y/sGmnHgurnn7A3iDm7mhnAFUwYxey4Efjm8yhFTj31rZiwzpCi
N4G1UnMPZxp6hJiSj1FcTKsEeL88jZEq3kqmza0G1X63aZF0tQlwxndswUuaPiNPkEQCGzXEwtRC
cNQzskK6dz9xD+H8f3S5af1cgIRwkZWNhS5OKmu5/ZUGpNLe8/ij6JETzBH3SRDsGekJVkSb5uuz
lkUb8KLbuKVDB38LwWD0+gkpxem2Z6wrn4FdEBPQ2Adzp4GrIPXEE69sNIJWo/CmMIFXznPkfr4k
7c/XVXe5IhbUUGm6nU2L32ljkUO9u63WFx/y8riEp5UQa4VV+n4xmgT1LhR98gLl7CB9/q5PUqeC
BEgsd11m3QH9r7DyF883I26CkeaE6YU5rozHYgQPclZICIewTCMoZAZ1TFEGbJgjq91f9NQDpUOc
6LcMCPcuWPd0xSMknWQb9hOGPGIYtOrRIbejwlI8jiaJx2aZ+p0CzLB5vn0oIt6DigizA8HV6ls2
6nr5DaLmD/H7n4ehD44g8+h1cm40NhjcfxTuYFSABiS/b6nLyjJ99duL3qKmHsiIT2VbOJCsNaN0
3yxYHF+Q7yvtY8dWl2Bn9e0uqcttwfeeDOSayDjvVkYomQypF49FtSaJKfVn5nZVGU6C+VCCuraJ
wtmPLoCEVUGvh4ZbSz2FRWfd+4FKv36qAnxRwOasV8oFcXWS7JAp0bxlOuTB2ih3d4W30+j9PHwf
csok47rzCJGrdjrXEfqc9nXZdUuWcQ9F4/SAIAEMXYsRMHwmIfrc79gw43+SGUg5ALjAtPXNbCFs
ZPjxebeN3UTbOUpHerGk1ToDWlFtPEy80UZ4+jmvr/njASZDt4xpgiYuSl4F8rhYOcYuooatUA1k
IUn0usM5YDixptcBeDUrfZiuskFL0yJnrYndoQBpgVoSeFP5/w6Aghh7ygB8aUXsJyj52MbVnNlZ
IcTeleyn9qOY8Y2AQ3nXhJU/n3g8xCnW5JywVX37VrT7OnE1tymWH4/8zDP+32aYB8VYQtylPmiY
gSsIk3WBfcsaaF4iRiLfWQCaOQgbQailHKL4ZGtS0Zra2JRd/EB9OrtuQcI1su0Kt9ItLz+gZhmN
Q35hATTtdb2C95OQkV/67ZsC0IBA6AslOuYS1+VQjQwUkxOcooVCF88l62GMsjUl9ajdslf9zoAw
Zch7fJQjY7EzXmb2ITk3crAL5iLj1AskCSaqyuQzFrwCk9WOOJAyHRMSmZK8X9xjjr26U/LO/ISr
IKl9tT5+Wx8pRVz6vx4xRUNhOuxC+JqJJ1szTXGDbstU9OoaBYVOOWC38ZSdisiBagWJExZFaMzt
u3AGGNvJvnoU1h2IAoEbMff4bZajUgyGp9nAObXR2bfsQD/3Ss1th1iFOm4Q6hQgEyLfMcZ27QRM
gPe0V3ziQGtnyN+jNBASGRfoGpKlIod4baQvAE1fIHSyEOP3A7bbAsKb+MQEDfR453i/XxAKCFEd
8qEjBD8jHP772EF4hVupKSuL1q5+3HBsQhr9p6yhlJZWkYfWXFb0B3ypfwiSNyuE9FF04jRGw8BE
fkU1wC3STtWGJW5KaAZi/rf8QhaOzWJI4kFinvCK0eRbuPHksqFaeLbByiJkBNlcFvEfz06u8ALx
7ET6gTWChgHBwJKScjfa9dtpqEWhIoGpznBtMpiNknU+1VSHfj3grngnLr8EulW+XuAhmJKBclxF
9MYCEPvfEaeS5jsflqwmiUEp9uH/7JMzhMtXFIZYC6IFjGI2sscBHExZ+Pi2DxUtet3mXKND7HYO
FBI/aJt0piz4B4yjYS6Pwfy/HPtKRGgwyj8H9irHSeawWqKCSVuFDUdY5Jp94t7JiTRneguv2/QK
roXR9TETlb+C8eVDPrL94P0gGUrQR6gz66PuTPVrWzfQ4Q6qMtosLJGSY70sb8peey1mDQXUgcB8
xGIQ3U8uueXX5iHs1lZBfktA3lYXrzSlHgVIeol7PGIOirle0uLj82ucUjI+GL+iWWqkqIeQ6kEf
WGwibP3mk+QMnoPzQjaScNT8ZHuAF7s+5vOk91OvhTt9n4cQa+nNS0k8mK+RhX4h78icz+Fr8/hB
S74LRLu12ZgeJKiwOzW0s2SXMPqz0eldGQs2fSSrw/9JefcG7ULSGwx7F53d5HnC6KL5H+ys+svw
F8L6QHVSO9hXypGVI97e3YtWHeMSSpa8mFesxMKZ4CNuYHxckDdgckIaNVJAx043Q9iZ6z/fqd3H
0VGBoGxAtqGWV29ZZUoXN0KlxZSOchXu3BmcjnVUNulI9B8jn708/lzDkYryEFk4K+kMv0Ot0vxK
55wRvaHGai1te98DkBVVVnJ/n6ib6/UzMlvtXKtkbgQz2bcXXXQRnfdT7MyxS7DO7IxJIops+LCj
ZmDaILMMl8EzdcjyylOoSozBcsdvmtEmEUdHaNJEWbCvWE9nmLyDEbDqxVdFGX3Dry1NXSXqs98u
DKjB3oPBNg5WFpagA+/VY+304ax+heEtnPM1ysW/nyO4yOhgWSGSyJCKgcHujZ3Q7Y/NkjLQ1ihm
/GxjpQkBlKv0+x+yl1JWwcb5ICLeZ+tYkl+5+Gt77D95d0GoI+G078MNsizZO5DS2vBREuzjyyom
+I+v9GSR/CtZK6QPNYVQrjw2GvBlm3vytOfSY/I1xReFT+/PAocBzNzwZRSMovOTXf/mIAFte1TD
wIHHZhgF77gZF9sO71uauulk+B6dRWztGoxQwHVXYy88z3PThTR8GQ+TLxVA/cD5zsb6YkM66bsG
2ffXO3Qu5AcwfmaeySejUHH1/f8I3kO1NyrjX/1lhHxNkQjv1T2DoeP2TYnG2WdFz2tct8ChdBXs
1155vT/sVEuog7hMecuD1Wf+KlNT6zVJcjYaCjgZXEh8QFGP1bfYzjXRpIejPfwO2Eb7izcylwDz
YgHPwCg5CMe47R/gmmWlnFqBkF4fqupeZgOBzvWOfM3xCMCuH8XZpStrti3IuQ9wwyxfq9xFWb8d
lxrYpBjkwCmYb9T5J+Qd/VvxvgTisoVCfOcqDnOxLn3WU1qhOkApAedMdmbnbrrN49UOOT54pdFS
7USdwz3TjZx90hEo8md1/N9d9bXLtu+wS9q4RzqRfiKEOufQIU9ttecBgc3lH1GTYHGMCDvxErR7
T+gBV4jWaHyJbw8376ZO5RCj9E6X+oeO82rcXMStAqt1JxKd+bVw8ZDJ+aompkv1fVK60qDsXNDZ
kMqVB6kJw/54aM5Yr43vTqk8JPum66QdmWnUJur0yv8m8DwRRDAb2FOCCoZMX5hi6TTFGIwSttKN
PCKGtNPJiXrh5OMrhU5dtGVb49CmSNwjoZZrnJAMLNoQU/6nHEZzgwqOJhKQX6dEkkonlLK9gy9V
oEjxo5mEFJTyx768vsGZvAvrM3tsVRpB4bPzFpIL30p5fM072Wg8xjLsV9Us6oEHWR/d8unWeQ7+
opuj2Jr8kbeWp+v8d1tai4Ctu0ChdP43t6WEqCxY+Q7JbuGbEPPpT5yN1P/tUc1tsfMZ0+JwcN25
bXUS2Q/wpL5Ja2PHtRBLCodB5NZrBTRY+WKGQTirAQKRh3EdGb31iSlOHrD4gABjtYSZi8DmmmXa
MOtxM3VbBLApLLjfcOBEIoHawBKm0Ts72Gqp2UhbXkihhWHKXkE1nbaTnEHNMV5Q7J3to7kx+a5Y
zzmhUp1xA/IzaMZc2IGeIzH3XNSZCarVJL3bWj+GMc+k2ByAg8FIHvRC9/gs5N3bK3m7PZMxu8hC
1NYrb+C9nQwVRfcUtw/s5QFApH7SxuE8EHrfJRsRK3BDAX+gdy/EcmshtBufgCLXUqNOLwGnTiC8
X1ETFkDgahDHU306UWbZ67CylQBrsXIC4juWdeXK6m5u479oMKtMdI1sq/D5AOe3HqWHFAgC7fpU
CctxX1jYJ0oCgw1ZGAtjJzn++L/0hQUzjjAVuWuAg8ZVw3tbqaDXfqLakXg08qGXj7Ykgh78wCUz
FhDUeqTa9BLZvvOt5KCy43Zvk/Le4QCU2qfhVLNg28zHodfWoDOrDxXmMOnSSvsNFKpnZ5Ex0/Kk
oY9lFeQsSPC9G2Ucb4HFWO+pi/aNSLxzIeJRF0FtVYXKul8pj3EHK5P8n8jNzrcpMAittDr8a//L
jOiORUA0613Gg7UFCZYdFnl6kRnKSIQLjK9csEQhA+YI2idIlpeytLh9ZvxF2sTkUf+Xs5P9amS8
DZfJfMmqv0nxZ2V/f5ie1VC9Xi7xNxR2mhFw9aWgNwEZmLR+jzRmFusD/zzh44rMYBNzkxjoSN5F
cz0WZIAPhBw6EdpxQSlhV8GG3xo7IZb6m9SGX5sdF2uLaA03oagpke40cXMkLd9RnVyYr8XsbLd2
/N8uVx+Xe2bTXWvypHivh60L/51Sx8Un0DbSEcRfQN7KmJruZQaqFKMIh+80SV7+dfjhE+ZkbI2Q
JyFThl8FiF9Mm4GbsfT3h647Gj5dPdYoy1XM6PC4K19LHQYT6hUldlIX73jnAmi2F4QjsM0ygtd+
LpLA3XVwrn20mUrGqD4N7U2Meam6/1qCKUE4ejTd7dJZoJe4SH4di0XWKJ7Lzw20itzGxiyV3NIc
tv5MQC3W9a1R/tjPrTd4h8gyuTqdDAs/sXWKr96WSlMdG1cMbXqX+MP4sfF6u+kqU+mbZ3DFDfSC
0szDwSUYfEB+hCbkatP4Y4hfWR9CvPwC3ylxVIviTVTOgA0Ix8sNCBNdwxRDMmoMZBniNIAl27CC
2Um0C2LxQzZxCK0464DvUJKDrMWD3+/WEHiwgfSGkfFIef/4nO3Vw5stTeEMOrPX7WNwKVAKgStz
wzQJNiHNfg1QlwTqvVg2DNtHf2m+nwKYMZz0Fs9cEsKuD1hYTm22/sQuThCZq8QfYqvsMvuTQBQR
rem5jgaOOmGwCQjlhPuIocWas1f9UxU4I8q7+HUTRlGpScfB3K0MMCRzFIi2lEH4d04XDW0l6V6y
nfuPNbkUaZxKNXR9bJlrce1jkIH3/KUOJmUdVSTOWSkDRkNNVL77EBfSnzLwKmqLrML9D2mAv+mR
3mhFdUNlSMHOsAvv+WaEmR36QR+iIZy21ju2IjFw/yrBtXasDMN0XlDAfV2hxoTgIEgDNRkAWVpN
3gpyBhGQMccrZiTd8bozxZr/vIuwJoANuhH4C2ObBhIk/330s93mOjbaK/19kTAAYP48cmq5o4xp
uxp0s6uT9vCufCq5xMw0BylRvEyrZ+/W4Gws44bpJvWuRDFPPNVqSPZQW0cyJ4RZ1EpUUxzOZI1K
O2/QPNvII9DI9XWa170n75N5ANVlgSPy70PNleZfwDkUCZhsOq4vYiGK2mffWccgnqkOJ+5Ao1LY
l5RhvA5ttWsJLRjHIlfAb/1kh0eBIguQa7ynKFXcxAsj11J2cmg3J7f9a31qIKbtZ8oi+DZ/YzZD
LBCYaPiDIw8LSjD7CTpbec+z7fpJJfo1HM6fc0qNplNgcKLXsZI8S5gQGRPJ1qO5tRZQaxPKcZAk
DitZWCytMlT0L8B/sbypIa2QAkxCq1oXLCzlHQ95rlcjwnwPVRxZ04TTuGYiYp1O5YmXFXWpMyBS
WJJo3uQ7vbD89RR+H3bRbQEqOp5eqf3+rg7pHg1lJUcuPjPKvdbHtlWqbukr/N+Q12CRKe7LcgTW
6p5yzwGked84OQ4UTlNPv8jih7MujBxXgstMxLjKCQyomozC3E9dXlv9CVI162PQTICfQhy9gaIi
OT6+GRhPTy9zRbdVWrEvn1Up39Glk30yaGOfXoxxCSj2WP9GJ4lZn9TcjWEJQy/JhRCjqWBLs0b0
6JV7wM94AzcjZN+zheIvuui9Ym5m5QFTVXZbJKEYeiG4XXnZh6IfllW9+A+KGjdQz6kYKbkrz4iC
F8zfTiNtnu/ZzFPdUyMgf4AjnCV/e6dvISeG5BLot6n7/s5qVMbJIs3WCTL7hQJilq/Hyc99HDxj
meJE+hqbQt6LkGGmOsn/KW61zKZgaklDXkqsy5Ou/iXrpaN9XKzauXZ2Px7ovTqCXYPp5KwRyFtE
0wSsZI6Kra6/rtpXL2WzJLKYzj7RqZX87fBcoK9bnAXn+2GhTjmoyfjXs9nLaK4+Y+cyxqHqdkYn
AyeHjc9Vt/RSunD47BSRzORuM5iX0TQ+Z98jE92YRqJXyaCrTV0jEe6nooQm09ELiYZzGCgdHfqc
f2PyrKkXopXjn+rABYb1T2YgBymMLRIF/Cjj3RbEAUP5vDEMhZjOG9veOxItGHTsBWp8zEX9IAdh
WT2KHn5S8fk5r36lVMYUCX82s8CODAdRQZub8rS4PqQ5bsh4hj4Nxm1ZQcgKFhBd2RzYxwr5CNuX
9i5UtErmu8sGSW7/RzE9l3fIPjow10j4AFe+WWHzTmqBdjtIn1beCcqLoDoaytzG81jEILqRE+qO
vYiE8PRUEnKZ4HZ1kJcDD0H1AJ6AHF+bRSnPUA9SNCFKUTO6icKELLZHAZuz6wML6Y+gmEnpJQ7R
4Kn7X3YAqc1/oVf3koRZrfJ2uGYXux5EgZOLsj0GA6UjtzG8aqoF3650uCi3d7rA9mETUFw/iDa7
EUx/VfDS8gabTvwsovODcgMyepaSUbQJrHwq9gD2FkYgrIJsietD52bdofzQ46+WxCB0OKOVKPnG
eE1aozTG3OMCODLeGer5a6miHJigajiCGv560zdBOMPsCo3bkXr5tqWh7csMlv/JwOp9JHX6/2M8
Awn83VqE6DCkP746iG8YP0QxKeZsazjJKKGxF2PwZiDq+5zpG+7pXCSmkvxV3WYfq7E0kPTsTJdr
fbBz+WTJEhijs987hb8DwqWc0MtKMx6t9K8F3Q8xmOE2U0CDP5sc9drgWpWQod9z0BNFS+TBa1BP
U9P15CTRyrMSRuB6WBtijY/tLHjhESPxDj1qrcKDrClRQVcyxKn9zCpzmKRjtGup8Q31hx96/fKD
HGD/VAhK8WI1XqSpazFOGW/3srvObYMGWfYi4BLTtRhUvXs+eRfFp1FEoERlGvDtUDdrFZKzV0y/
zf2vmbqu2eA+8uQQFvr8YYpQ7l7W5tVN2SwW6oZ763U/QrXWmwcMiMtYFcQqKoA3xkd8u1kijHEE
CyFvcebiYyV2grlQCmuTmwRcfUVY9PBiKbMOuGY1IDH7gpReDZe8A/UOLb9r3VBoG0TXQTXLBzp7
JWd5SwKPSij7xxPhglazw3iUXS8VSpU/iFVZJnute3GCcJDWkM4rymEl7A5gHXeS2seKgfcm44iK
xKkF1rT/asMriidev1oKBSYgj4HZckaee8bJ3Plk2Gq9i9RVPiW+lgKQ6dsjHXKN9YyXvBHhR7lg
YyzHhSlicnhNFYjYyhIxbTxPxreDJ568O0vvUmQI30s7KrGS0NZaW8MYRkQQcfBoXTNatSXyPkcJ
dupoQIeQb/3vqEqRpsAaPt4lL858Yw/+lYcSEHLZrmbmUtXfgGIKkFRml1fY8YnseG3g3PeHboL1
NO2CpqwhpoFYixX4AUhHM5K0powBEtxhYmjwTj82KpvL9i/ghibOPiLGWx75Ginkr/WlMs15Yez3
7BvY+iu0iUI6GUqkmxBd4zraSdEk40fl+YWvjruGyGOevkCeP6/V8JlIpCO22tZrSsGO4Z6aT78N
dA5SXNOHTqDrF77cTHIC5Dgm7LLhEeRaWUO/AjfbrIqHhAiFGIK3jQxsCugvMK7dVCIIzvkxce5U
m8CT1JD5O7T7a2xE+5QONS8+414O5dSIh8AYVxa2hRxosKbd7ISF5dx+ZkEHYxnvWvHteQ3TPZW2
bv/gHLUUVlIHErERvM7mdqKP6LmfoZKNuu9bUUPDTvaqC6g8MFke16jzH+FD07+Ih9rzQPunHzmk
nm5nWVA7Sp/15Aaquqxdw03N61fW5Qr/PQU3512FCK/Foht+d+8uWQagxrcfL+vlf/0od8Ms2p9H
s5gBySaGfFFk7LQfa1cyKYdFKBsOWvDEivVtJezCWhYfzKB8fEZELYHhAZOHf+hOL+crnsmVoN1f
pBjCFVm5Rn/j6HdMIzCjMFXHZMrvjvTy5Kt2qzDVYEwmTOKKgkgIYobjRRPfmn4O71GNAZ62h+Kt
yq7rUOCnbf/wp7VuXlYGbfvOR2ppLs4UEibs4KLU2dWOqeWuMM6VCmv96zegFU2nCldgBlNGeShm
xQ0XBVXJ5xpGyiegYdEaTYq/F/yH1o89XwlT1ROClD7CWV4CqWg3fDPEVCqn9g7k0n1wb9LZ7IG5
vbw8OES3OL7xx2K6keIjy5AQ4nhMMQ42L8F7ZZKB9Ggw48+RndcnWcMXfPj+M5rZIpZ8LPoTYGqR
zBCnjsOlKm6HCkG9MNFjpD5hLfM+Zrai4A2B3ulL2PSsABZ4X9PmUmOU/9ogDFR8AYix9bWJdA8K
U9x1ENfPPz0nrt+GKp05s0zd+h6YgnoCFo7kbw+j3i/dTMS+97InarT2q2CXv7gqkC2ehdv33Att
Rknd7jzffaSmzZHJsva5Hql7DeWWg3Mo8AObQI7VmWgRVTtcaAP1xHHcsrkvQ/JrYHjZCI3ksl8c
gmqaQBV9k+GW51ArSxtq0tUhU5v036qu6Ct7CEW0TkMo5XJ+ZoCesqnDpClDByaCaSIuSAKGuxsk
2wACzD3vVXi/KLXW9vHW4yU4D1v7VHVLQmWTN8qwHCxdtirmNU2ux57kHgtBDfzMs29vIETiR0Vg
/XcISzuTuRasb9jjxljevubcVa4HNFzKL/Xs5KuThmnmcP+vC7AlI5pwGHw1IsJrqB9JJk/rLqEM
jZ1KiE/wMFboIVU5ZnUbtsTQTPCj7f/EABD6xSduSvYJKHCIguss3ckaNXUoc7ceb7o2Sq2ThltB
Sea2lVUothJO6nhGPpa5nWSZmK4HiPoU1RqoIJ/UPeYHMfOZ4aAF6fi6YkyEn+kup2KpYvE0Y+rg
fURt6/hc3fAN0odQOjRKoLimk2+pTLBuwzhOamHzVuho4zrh/enVs22xmYNq/+GI6LpVIcBpUpuy
YfQCceztpNEX1M/3HnsO+lFPstzZWxkDF+QnMxdDrN30EsbV4o67V9AIMbV2ZUEDapFzzygy700H
D3FKXQ5wK8Ymi0B4sbKpS/AK3SNChnpK2q5WC0MirXX2sdrhbieSDmllgKWqst1Ss7VRi/gRN7ei
Wf2S1kV5H68lTjYfjHyYpWZX2nq1tbO/x8l4007vwQmQxZ2xKMn0SwfHVX21ksmViEerUpt52dgT
IIUJSJPbov5h3LMFEkWUqEc1PvmAFKGOaKDuh+VQTpbORiMyltT+5/WdeNoZmgim1SiGTyZ9a35q
85PIYVl1wui6AJHgIN0gNw6piEm9ZIb48B+Xwr/ds5ecq7HM2YcNUnhgqWVT+/vcBUOdoHrJkza4
t2Oa6UhPAXtss5XLK0aNwMbCb7YszoWCi4uCYtqu7L6wgFT8uMNciuXeyt/AO4Dz7FRNysLq5jLv
Lzk2QxiKd9IvjIhJ92fJYZpBAQvwfuKZ5ySaHSfLXaSLxiRSMTaGUe/AHAGsEX5pyxtrwN7MBRhr
DFImTR932A4UWN1KgSZ/eMCI/IQ7r/GsiVSB7rnNxpp2kFgpTHLWOkUtEB4N0JihYHYtkh2yZ9gm
no0n/X2ZcCzpg0RTiGbM85KQ2V7JMSIRBYz1ibuqh7tLPntj7+nUwdAYBRACjUim/Srf0H+u6eUw
mAy7cSV2HtJOEg6KbDg2oriLuJsSiNeEjPiktU9yWM/+0HNNot2kgPHE0ESF2YRjTdjcD1HDDwYn
mU4zwvMsA6tI+sWanUPzry4V42xxWx1GdhvsRmAApDArGuauFKCOHY6ulglffoiTxNIbtIEH7avw
WLXdHOl07naMlSDe2d5qqLQLUWeZ2141+BTI7noiaATDGHlOeYUZZXKWCG9GiZrlYcRhyVr3lDDr
jGMbSHGusfA0Z9eWAIRrGtZsxnU7qaqbDRTw3uNsrqjxy0x+R0emjYeHsA8rN+xKbTEnw/4nf42P
488B4rpvC8vhiUy5zS3C432Td9UsNy4mwXDDVqHzSJtMTAIHUGbuHufXY6CxgTliWqzT+FVcJdKX
wIvswnMKLYsGj8hyyTbWeS25XpLshfEvXjrRKH585SlEkOqiDz6r5vvZCj5HPlx0T9OhkndPtNCW
6Tqubm5JRpwAGh8MLqeJ2i2RlUntcMt4T0jjQ+Gkp/PqZR4Y0/xorWxHQ1zyjNvflAR7/iHLYhGw
wKIBjSAmmuK22yHd/78UEGqpU84/60KxSJCrfUUzAmpGjqgxli7PgjLhuIgX4kVfoY59xjMXhXr4
XF8FQGLAfAreN5Y1Myikn/FG+BKA0zlrgwNsHDMBXWiRFkoavZjoX1+tDf6Hpnj52yJyf5e82qrX
wwq2+/B5AOJ9DaAHRSG4m3X+pj8N3qyiaVC5PQkmANElfNSJ9OlgTtddSj3LMQbjY66RKCrHBuMD
uR71LbSxV889i3JSekV9eaOJaWCpo/JwE5/OxA/L68xV8UCwL+h5XdRQNS4tnkChNTTN/HNkvtut
0gRYuL+axaWReedXP0j26wtqNKwIDRRzYhqq8UF/STTbeCbB18VaEgtGyxXPgh8yx6t2xvfL1Ms5
7sa5QhpH0FkEbb9wemy7lp/WXbHAnit5WcdhKg4h76ryyq/fl0Bb8Zlkhfxu9zrxLSa6tHWWMrc7
CukHa7iWFTSitbEixbOXk3kYyc+T4HMlL5kfC6xeKbbj/vmquLyivL+2AVJObMsGC1yirfEvnGIc
BC1J2NkEYGA1M9jSeJm7R9ZL8kBr1OCxQriW0gBfqLVQFPV4Dh12GZxd/81AgYO8m7uuNaD3H/3W
WQCWAekheWNf3lL+g39nUADeCFwlXa+nr2zp6wxRNQEoXm4rwEZVzZr5LjxSr5m3LJa+1dkFFur3
nhzRl1e6zwk6QITJHhar4DLs8og6NsCT/qYtNuAmSCMU/pgLOF4rK/FiFEUvjSLtKCMzDpRMTyLe
XHAladSfrN2RmFVEieN4PuEBTanojsNL31Z+RctWs3tt3H7AfAKZdaqdR5UptVqNfh6IonWQ2IcG
KXi5jC7wRxc9sTQxxXBv0cUJdz+f2BiU4ewnW60kpYf+7meFkLhsnMKs2W7KvGAf5IwSEkvvQRhX
oW/UolXM03J5PyQqzQ7oCHZPxjkREmHGg/mkq6Yz4muzm9GfFkRwPyWbk4hEkfIwGOpJgB5qIcq3
zt25spLbn4ITsoj8lO0QsXNFmQaXa5P9o5ION1ysflrPhw4hiaL0ZzTM6e3ghO7HlWoQ8mGgPnjH
7Qtszv2LvPGsEfIbjiTmLvs1x7h13v8vyy6b+hrzc+04QKyUPBXcQ3DGOiz3zFzTp8oXScSSTGdA
xTsDIhUMooL689IOkuUu+JvKXUMfv+UGVZu9triHlTR5tDGZ+jVq9E6GX57I8n2MMEG1GKo+dIb/
Wdt5c2Yfgpg5xcRMYf58+HtQtoE32BsI8rM/jbcfP/hqgt0DUmBkirZIvKocKn2XojZ/beQpyDoh
VDUghmZLpZYwz1lIIPcS6EFIk/svgQRfDuiWNhzjaEetrqczGEPZYsAyArhT7L9pX/yFsReDdOke
eKdg/TujHCJLuoniF+ocrpBsYEKZnqTz+aShxctEOOaWB6oxK5wHs1fYcBSnejh/mfUhFPVdXj3i
kE/I02w/pkLgrqUYIRljbEIT3eAGEQrKXTHb5+Mi933xWk4hclJ7XwLFXXWiK+7FCy2Ud+XCuvUI
b9FVCuuQQxBAxzEojshGTGuZFKmkGQY=
`pragma protect end_protected
