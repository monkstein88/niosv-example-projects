��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a�����/�	v�+����@ɧ-3�����Iz�t�܀Le'H>	6"�U{��9�bEɤ6-�!�V��s� ���m�|����~μn���}�iԹ*VC�4���m7���-� �7�o�d�0w1 �⹺�)=k�:+5:� _M�e�$�"��O��0U̅�iZ��x�K�~̏*���;��R+X�="+$Y~�ml���n�H���K1,���0�ϔ���憲e'oN��D_lxY��^PZ�#�C�e��Au�֝��2ɤZ2���ܵ� �o���ǣߜM0ځr5r`D.ɩ�
e���
�Dc�����gC�8$����lc'�'@��A��Se��J�oY�\�?f�ᕭ�o0�\�O��H�$���m���M2�M��J��?�c��ˈA���~=ɮ�����D���B�p��;�e㹽yU4-����_8����p�R�C7�H��;v��F��5	��zMV�I�xB�cȀ�j��� l�{�I�e>;�IT�NF.v2���hb�]%fzy�0���#�%�GNאsXU�թ���*��j�5x
�P2V�?��9}��=�->���x�/#v��_�����J�N�(��x�USy��i7�4��J�ÞQb���u����V��i/��R�	J�,W��r����tx�E�r}ӣ��בrl��P=��������1+�&r�W]�#'`��5]h�?�G�i��:b�P�Ǎ�;�׈6����r�R�����
m;��V�j�w��^Q�Z1�d�p#��`�h� ����Ҹ"���'�1��o�}��d_��0�^$-9S������b�I'Ѿ(==� �����N^X39޻f�z�M߶�>m�84�G�d�|6� >��2'[�a[g� �oL�(Y�h/G���ܚ�ղy)a���l��� �d�,�f5�gFS4|�M8l> �����0<O`q�`�U�X�$.?@�S�xm���h*#���_��)��a��i��<g��Mە�����3xt�F�����ef̌�����:Pn�� EM�é�=����/�̣S1��$��<a��\u�!/�\����փ ���:�u���־��Q��2�sƴF�X�������)|=ZϠI�2É3�K�%3ń��q�؍o* t"it`�+��7��܌�G\{�ף�O���Y���}9:\x:��8'm�"�W>@����--3v��m�|�6P�yF+�O8ە+O��&XV+�������I^Q��C���)X�1���Wש��d�Am@!v�4M2P��=k�	�S!�٪��PP6֒� �l���u����+�#ϟ���P�̗(9�@a��9�I�N��4�vX���S���R�F�l���P�[����=#Or���$Ӏ��������l� �mfy��_�͹�e8\�HW�5/vmV�����.�9�1��,4p3t�&�5�q����˼�y�U0�0!)�Il\���[���VE8�����:G
�LT�)��{0�<�5 L��f`�8Vΰ
Un�]Iq���& ��[\1�!�B�������V��A�J%�X�KvO<큌}^#���P�^�(&�C��0v���l����7�{]�|&'K�}��aU�N� ԍC��vц��WZx-;��'������mG�m�:��I�<�\�|���$^�# �jCI� 7�za�$�ļ:r��L�D����%�߰�
�1����O_�������9��)#���l�5J4$u�\�0]F�UҶP�~����c���̬z:j�4թ �� �ꉺ<b9Ub���I&��S�R���o5�`K�,;��	�fs���^7����]N�ʘ��~.Q�''�s�����W�'K�f����k$$�����z���f,@��)��,����y<�7]��_�����z�?��L��q���+`�:�զ��Q�޻��gk�[@A?��s���� NrD�[�8���6�DidXU��t*`���%!�ZR��n�O�Xj�q7cru꜀c��3& k�׍����˨i3���T�S�������p.��x�b�tc�D~ZjX�j�Y��C(��}ӡ��,��<��7h� 9����E~�^���)��!m���򏉜*Ha��m��!rV�1���r5�Z�R;�X�bV+zA;�s�Q����'�r�Wбf%g��9`�]��p�S����,��أ�����٭�}�o��v�>���i����?5T}$��ޒi�׸�*��NZ&��Wj̰�x�nS�:��G{��^|�%��nV�Xs$��!��N:*�x<�ΛM��m����P�E�Ѻ4h·{Xo�8��2vݞ�Xƴ��^|�}sf;��:$3jyV6;�(�U��R��d	�4��.i)>�o��	��N
.����w�H)��y��'-%<[nq�U�o��Qs���(����8�c�[t���oyh��g0�fJ�x�ܪ�f�H`Ug�B�T�����̿A�-�{�nd�U�h"�C��*��Ϗz�?�("�qA/��l䚎���ȯL��t�pFr�=	�4����d��.��憺�m�ݷ;�=�MD��%�)T�Ы0�*\���:��=~)�ujH�\�{GSlXd�����vv	���CdXC�5%op�}*�e����_f���(sEQ� w�]�%XZ�`��\�&�2Ș��GM"���'��M0[lk'��r��)���n9���P��$O�o��j�BNf�9v�&F�SO��W�*�g�wV!$�E�Xy���<9zÍH΃"Q��:���ڥ=:��o�;���>"Lt��Pv��O���E"������y�cï��kE7TL=��B=s�N�@�4�(�R���vС(pמ#hR��$-�d��f?�GD�1���|� ���ly���ө�]��}�;q*�\[�����cEv�u�5x��wG�m
!?fǎֺl�>��ס��l��zb�M��0����۶=�{�TT��z��]`��v^ݏ����ыm]r�O��&NyϠUbpJzS�����I��8 Z��P�Wtd��t�#h���
~��,����\���c��t�7c��3+!*��B��0�h������8�`�����6b���d�F���qV�Vj�!�Yo��)�A-rR�ϔ�w�{^��֙����q*y�� �A�Q��&e[���	gJ�U�_�%+�Vl�
���ʹ��nÐ�_M��3�帎�WZ��XUm(��B�}��|'�w*��Hz�}��jdƲ�����2W�~�^�>�@1[w����Nƿ��4~����s8QD.���|pwx-��I�=���g��
Z
�6e�!��wk�:+R�]�e3��ߕ�wr�<?�͖^�m1���D��?����j��V��?9d��������@~�'wVt0`��͗��@�Og��3�M�Qׇp�$02b�-��_0wv��F�)؄ϫ����%�K��]M�N{E����3b��j����5���� ��ˁd=��щ��8��n�<O�f�F��~#Eh4|��'\�]�
�8�^K�����{�m���X����ɉiy��t�b�C�+"|]�^ȾK�;b��A����V�η,: uÿ�iķCq����)�Co];���{�9�K��9��.�Ou��X�5\�\:��i/���X�-=q�r�D��=�0�y����w��r���s�0�~l����}��/άS��0/��i��T~y���H�e�/{�������_���\B��z�{׀'�k�&��Eͱ X�!�5�}=�6ܖ"�0B�A�r@�9j�+I���%hA�"δh^�H�:[��&���є�c�0Z��s����@E6b͂y<���c�V�wV��s�"^L��n�0#4�d�a�*&U?��ozbGO+�y�B�>��ki3�Up/NЗ��Q�X���z��A��� ���{u�+��Ć�r���&jyA,����_x���Sy�5�q�b�4'���Ď}��`@����@ R5�Z�>/.�8��C�Kϒ���=��ׯ��Kmh�y�z��"��W� ���w�#Q���c�=r���p7�~���V����Te��U�t����-q��Pw����G��/O�N������1"y�
�{�vi�e����*��t�y��=[O��S b�[������R`�j���܂���
�M��l(�Ԛ�BH}/3gq�@��,=!��/O��������&]������-j�W߆�dC�%)ᩊ��Ov����5>�s�����v�T���
a���i����̈́[60�Jp���"�g�#�%����zP�U^c8~tPP^� &l���T�K@}���n�*�M���T��u�&i��	&Vy��������Ȅt���v��̋A�zB����hُ|G�,ə(��&�^-C���R�\��^z�t�0:-ޖ����8Ϯ�{�$�qi�H��� ��>.�P,���w��C+�P�4�+�բ<�����6����B�ط��R�&ш���m�r:�ϼ9���:\�.����s�OLÅ
��Ǟ�,6c�9���\���Eы;r!�����۪�&�+؅�_:L��9۶_餔^Vi��������G(����(��U��KB5�K��(��-u+�xZ=�Iv(Ba1����D�����I�Ҹ}�]W���CRnr��Wv@k%Rr1},��̈́6h��o�� {5�l�]�eQ΀&��9d;ԩ��MQ�j���I	���l�v] [}$p6��K�Z��mZ�*�Yԉy�B:��y؀��X�:5��B��,�|��gcԊ������)�N�q/�[� S���s.�'`���1�m�F�pI�ҧ7���yi��y��P�<�~E	$�ڭ��{�EsN7P�;�f]	�%�r�%�1�d�;����PMs��qd_�|��[�Σ;$A�9}�.95S�;�)T�PE��3��	T#�2��j�1��0_�8닐���`�sL��TO�Uێ �QK�Ȋ�!��5��������^� dO�"#`���&J]�`��g9_��Q�y�!��q����N֘�Jx�/R,��J6F��7���/�'TITG�����j��TϿ��2j�P SC)���g#���%Hc;_v[GX$���)ώ����R'�\3���-��ԓg@6�p���`e�ԩ13Wjsn�|*ݘ�T�-d�J��&@��é��d;���ԍL��Xx��x��zL\wuKoJ��2��@ �w"�Gl^ր�c�ћ�Z�iI��T���v�+!!8u����n/���R���k'2tz�oh���>دe�g�
!:�+C��Ju�N)ZJ�z�É/������{������Y�=b�RNq�!���	�PHt�?������q Ϙ�x兠3H�=3}�A|u�}�
_�l^*Q�(�x�j%%��@ ���.r���J��K�`�d(��79������/4lP�	�z�q��jL�jٛ�%�:�s�<5��I��Q�%�zɻI�Bs"��%�"�±t�.'�Ժ�1�O��[JrL$�����E ~FK3�P���WP�6��B�D(P�u��R��&�Ȯ�8������/��YP��*4�S"���`��N�7��֟J���	}������ N�f.��TsN�8�"_{�%.�~Q���҆�2�[��	�9���W����j��0�|���w">���H#�����>�Eg�r_������Y����d�ˍ{�!��1P0�v�\��T�mۢC7��,�Y��4.V1Ӊ�Q7�SzqI��XK��8����w�엥5Wfv��\�M����{/��<�G��CϗN�Ֆ:��A#�8<�����
�pf�c�����,�2lO�E�9D�m�7�. ��.��X�.�����;+�&GT����F���S��ո�5�>;�zr�]O���D� � DN=z/�?�G��O���Zv���iJ��p@y��j�-\���o�lt��w��b�\��,7F=hsP��o�(���R�a@}N)�BNisd��g:7`-[*��k�ث1G���:�:4��!~�\�,l��lL�cp`J�ݴ���L��\[.����`
!Ԡ�`:��HA����
U��{pxV�<�&�/����3���Z��р�Ǡ�Dh���t�f��k�meZ�%������Y�Fh������U�<$a	�� &`^ê�����h�:<=��������j���aA:H�.L{��|A�6iZoF���M~\�DA�y<�2ѧLֳ�lB��q'RϨ���KH�{P�n���e�p�/l�����[@ۦY�Sbv稶��Xƕ��ٜ��l?�<V�N4���⅛n�i�J�r���E#����򸚾�0�����ˈ��ъ��ȮY8����K���]�Ƕ �������%̻�8w�4������Jsz�����g�*Ƞ9�I�0�w�m�c}�$��Q���s�d��U�� ���J�g��Tf�+�Ս��@��r�F��F�A��L}B6 �(#,�t��>4�j>nx���֭FV�F��n�	��Wx�ȁf|�߇NGd�\����.|�);$��jSg�+�L�P�sd��=�f6gɧ�T%�4W(��i�7֧��k��=���Z�Ε�i� &��A���|�`�XA��;�5^��P")�(��n���`!���ؙ���dԞnC��Q�A�y�����o�P��N�[�P�D�?�(�P���u�`DPWto��:�K2r�*�Wִ%�Nq���Y����&����s�J��><�Z�Y#p�>	�Y�Q,\5��I�,�s��ڱl]a��K��6q���@&ىd@:�/���\9�,�Q*�RX��۫-�.e0a���G$���a��ur��4n����%�
���%���k����y�%T��8��N��`3�y�o�8\�h�R���}hO������+`�מ�延�z/\<�z��-��*��|��Ԑ��&���Oy��jM�~W� ��OE>bݎѧ�c�T�p������>͜�@�#�f���:���p�n�.ۭ���'�o�W&��D�9��N��DBS��5S��$� ThL���:mb��n(8����i@l�H���p��0)ԭ����v�$�LnfCv8ۂ�H�j2a(j��>j����*�S��v�wrch�//.�(�1�N$:H>aB�m���KB�&�%�v�Ě#?����A&Mg��bu��LDݓS}i�����cB{�|#�P��o���ȜVI�r}����ҀT͞v޴��JE��
�����7I�p��W����\�y����JBx��������ۜ�o����0g��	5�r�����@4#zD�b���O�07A�U)Ȃ��4�vU�QJ�)��M����(`�g[�W�[{n��}�p�L;V���F��{�T`��Bt6+:64�jY�8DK8D(d��%96+���:A~WQF��@�J!�F]��C�xm��|���$������-l̇��r��Q��B�z
�'�K�oH��_�8�W9��k��ˤ̓$��i���u�����0;���#QCMA��k/�.!>e�P	��`�f����=�7��a@.�*+�\��S�l�GQ��,Յ☝�L.��l��f�T�m�քB=�Ξ�l@�@}��Y�(Y��L�a�e:�L����$��,��V-:Xm}CV�Q�~��u%�Od�&�JZT��{�����Aݐ�h�t]᧞Cn�\�@���4`,���_w�#bAu"̵���']��b��(R�9�{�	$��`D��e�0���w�$t\�O�𑼂Cqi#[�8�ժ\��(,���+ǵ$T��Y�*�Q��v-��3�L?�_rv@��Gd��O
�Rw knr$�!�=��J�'�>z�L��K�76��1�y�>9׭���`6��Zh$����J�D�Ŗ?�>";�_�Վ.h'ж]������U��sp���1�MT(����}�T�~���ЄӗC�a"�7Wj���ܻ��*���v{�5���Q�ʂ���+�al��i�FR���6�w���̙�]���.�,��P���W�g��\��a���0X�W/4��*[���8iֺ��|3ŮF���T�~�Ȗ��uQm�h9̺B][���L턣�}yLn��#���M{[��*9I� v^X,�p�����`T�R��/�J/����X���d� �����9�]�Ɔ #����N�bė�
=Jnq�fAnZ6i)����Q|t�7h�~;;["�,ȸR:N�.H'z>s���]>v�B�T�ϾÒ�^LQ,��{��	<<Ȑ�<���!�P©h!���t�����\�7��u����n~�8����u�C�2��P)i�]Wt5����=Zx5k�Z�<��[`j1܋y�7a���G�>SVy�R5U��~�:� �a�3��e\<����T���+���M~:"1�{���)�+QR���6�v�ii���]|I��9$m�dV"�Т��H�aM�쇜b5�@����4.F��ۗ<���܌�.�H�x��ur���]{���`�^t�A�vO	�����������Mv9�l:i6� ��(|���5Z�ņa.qG�
���k_ϩ�p`�������Q�J��D��ZC�d��W��OX�ڱ�y��m�-n��f d�zJ=-	�r,����9����qU�*��7h��9k��$d2�rW�曡�=�m�`��6҆���f��r:�����W���ü�/IK0�����EUR�"M��6{�B/N����(��%%P�%b�P��~��y"3�r�i�@K|�b���s�s���f��UI#��yaQ���z�����=i�y�R ��H��v�|�ۡ8գ�m�}蝎�tXZ�IS���1�34:��R^_p��3bn�w'K�Gٕv��:t�W�B�I�~���,j�Ue"�d�kѽ� L�:�^rU���=�q�W�ƺ�ʒ�GW����y	J1g��JqO��ƙ����ʬ�š�9'f����(�T�8�K?������Nn�	x)�,ȚI�w�Um���o��8("����0��Tm)_�����t�ͼ-3����Z�B�Aw�ҫE�q���1��c��-&�]��hl�zr�82&�~�̼a�{z��KϽˡ7c�s�!<"ǹ#��,k&�.�@��t�2�@.:����VŮƢ��_�X����6����n3�X�~C����N��8� 2�������;z�{?EՍmFp=C�3���@�9��}Pl����(�uɲ��ш(+�а��+���N�a��s�{�c��$�yiϸ^j��!�ۋ�:k�eU�?�q+P��"do��a�6��i"��S�C��������X�/���֫*���j]@��n��$�J��b�.��~�ߜs�?��A�.^σ�6련�T�@0mC�x�������1�Q�~���{o	o���zR��BݫφJ7�2�XŞ"�<�<QkJ��du!����D�����;g��C#ʕT_��W���nE�IZ�`�#�����e>��r�i�P�m�-3�G�w-[A��1�'5D����=�"���Hd�a�����(��G֋Ю5P���f�gQG�=0����B��3��H�����D�2t5N*��jw� U��z�1�T1mWEZ���)��8���kr���ձDa':�Ñ#]��x<�lyЬu�T��{[�Vr�%~G�2Of3� w�;�ݸ�O6)�5�w�� �� vl�D|$B|R��3�8�/2��oTҪ����g�Ce{���\8f��\��~$1��[gf�#<ڻ�����H6D���yrBq$����y~������;z�G�u�9l|S�A}�ܠR�U#*�u;�&��+3��?�mx!�t��ꂁ�<�,d#P/���	ู�A�H3V�����oȅ��1�Hg������E�U�=(kr�dzHA��j��u]�8CC 
-z:?p/��J�|�T�!�� �D�(A�$\su�<�gSɃEGĚ�]�m���S&�B�����t׾O�B�r�;���+Ik�1��RX
l"��g9@�\Jr7�W� �k�n�<��U6ޒ-88���n&��c'�c�Q���	�ˤ�=|��#Y�*PE���h^���>/���-����u�T��s0�¦Ge���7�ɽU������9����h�m1���ߨ�m*��(i�"����b��މ�
��������^ڀ��ED`�j)q��QSu�+�{�F�h��Ͱ��]\J3|�DH���9������D��`��w\2l����bat�����L�i^��w/A�Kvt|B�76JX>J�o!y�]5����ds�pqӆ;K�'0w�m6��TZ�V���$����*��s��p>&8}N��]>}�P�qIɮ�eJ��4ՙ�'�V�M�;|�m��h���Ҝ�htɮG�R���W�VAm:|�p�&�$�_�ȗhy�z���.���8b��C�����A�3~"��V��&�mbk�-�+�k�љ�{���@3<xX��u��C�pqȅ�+(�J,R��q����[O����x$��EiߣNL^��} wO ��N�*�i�DN�2bW����}�b7Owi��NWՒ@�E�]?rDHA��{������v����bF���c��{ ���X�[�n����P5�gz���R�V�����%��
V����NZ�K�Bku��o_�۠s��~�V��q�k�R���׬���R���x��(D��z�}<�P�D{Y��g�?`�%�˰<Ō&MT���Лo�D_�%���U�<K�M� P��Y�����D\�6����u4`j��j��Ŷ��u�S��n���po����s����Q��5Iå�W�,�0�ڃOT�j�u�����M�j}�a �J�$�E��[�~N�:D��E��dV
����m��I������V~��s�L�Qǔ�"��h�|��N.�j�캄��e�q�矨��[��x I�����%lE \_QJ�aer�k�-�6��,T��[�Riߙ[���p죝�i�s� ��b瀻�
,��X�~B
Gf�������9��g�Q���tf�+��E:'XJK�л���� ��8�ȨNX�<4>�R�츛�ZC�p���#����ƽ�/�Z����@��/�)}FLj�ߘ�%�n <_���~����ȌN>��/�ø�BJ��,'���1K���u�* b��E�(U��{'�����9��
�E	W��|�yᕙ8OF#ЭS��e�6E3M8Q�0�H�sJ��F�:˗&�r�J�-��dd�w��t��IcH�}Y�?�n��i���e�����y�n�=mVL��D��y��A�o�%ޙ��|����54}:���"a7%0&��u%�EZ}.���o�j���৏�geS�A��?j�:�U�a�)S�����ނc��5��~^���[�i;eu,' ���w�_�g�	ٮF�����	�E��ïkc��1��|}`ɞ���(E�u��:�ł���٪5 �k3����2�S��"�N�[j�;*V�t� aV�'� �Q���H0���ڌ�B!�kr�{d�mCCb�!v7���O�ħ�=��`�=\d�^~-6�_L2,5�PcQ����!Q���cS3*�.��#��@u�Ǚk����hI�vmA�U6��b�U6E�i�H�	�Z�p���U�q)]�f�g�;Rx|��+-̄^����b�67t:R�rH���gY~3���LhvR�M��� ��,����$D�ru��2�]�Ҽ�d��fL*��<U	�<��9��Vi��+�r0'��Ϥ1�yv"��m0B����ݮ�>�ve�����r�W�/�WO��c�(�X^I��h��xA\Y�m�C�0�A���N�?��ǁN�X���o�d�ԪOxf��Ӿ.�$B����P>�`ب2`X�v&A{�]�5�C�R��$?��8�v��w`t�s�x������A�"���Ĥ�m�;��H
�M�>Ѧ҉���f\��tuDchb�;���0M��p*��ʧFI��������뭈���0��õ��o�7��ѨyP�]
9FE���<$aOP��=�T��
2rI�jvz����FGY�͢a�K��hjK��#{��!�1�1�K���]i��i�Z�d'�j�UQb͛�O�Z��������beDn�1*�V�R.q�����-���<�e����3��.;�NB�².��֊7��-�է��%�J<���`X�C���oD5][=,��
��/�z3��c2��U�d��'��^\�����2X\z=��@�g�.1�� �(t�p��'��J�ѡ�mPG���`3�cT��g���pr��Ap�q���;�1���d�t�#o�-�
М,%:ƋdW��_�Gs�vuQ׻�0;��1b�W�]�PP�5m��]{�㢹,_Xn.��e�6�t����{X+���u�.S�Bie�
����1�vU��9T����׈F�������.�sF�M�S}�v�6������c������CզW>q��Hq��<�<1q���zϹQ��Ͻ�dq+�7C�Fw�ʣ�d�Zr=�[���쥤Z���v�>�?�a�8��s�������1�}��O�T��M�J?S�z�^���%Tf�E��hH30��85�����?Ny}�NIɛ_EF
0��9��L�[�L"͍�>�;���֑h�z�e|�� �x���M����cۚ����Qa�2�I%g��?x����G<�}%P�������,�����6M�����5=�sIFi��K���7/��g �SY�#���aG�i����/Ǳ�rE��� ̺�I�?.���/�K�����f��A��,�����{g�r��?� ̀��.�����CKi�ˍ��q����\��:+�@�-=d�����R,�'�0��p_���/�㈢�kҷ�b`4������8/?l�mO�L�\��e� ��W+_?��Vv?��T#���A�6��s�#МE��S������I�UT��ΐ\� tHn�h����+�R�i&��|���^FY�R�^��ւ�A��	�A����9x���͖͝4���� �n�gd~�0�;`���ɔaD�2ލj��ߕ��0�\X����V�"��`)���O�KcrbH�cN7O(��v����ʣ�>2�8'ɕ02=��k2�^n.��<�̄�$F�E�,�6�j����j�Q�F���Ό䴚�L��a�ݠp`�<%��5�`c"?�'=!�\O�E����?/������^4(�+�8[q�i�����)�&*�ّ���h��2�e�������Ғ�!>����š�-���9Ϙ1���d:�w�$�P� �t.e0�x�K�#-�1�2~;�������*�s�Q@G^?sj;�UIk�o��s���9Ga%��-w��
��3²�O�	���o��z����V2f���d�$Ō��-
��%�OX����L�@�㴟O蛧��d%� E{J��
�5����{�.m�y��!U�d�&0� ����Q6?��?V#t�Һƣ�Ա�Gq�,�����]K�n�3������0x=�b��?��XL$��!_�V(w4F�L)�����.�<k��O7������Q^�Mx���ו*����^=�9�-�B.��g�0.}2^65���B�?3�5�)��OF�<�S+�2`�g�K��T��)��4&�<[']���+���ңex�d>�q�Z1���97�tD��|n��t&�����2�-
���|c��?�\7�*|����n�v�nr�jzH��zQ�(��n��D5����SFN�|�$R�Ԫz���L_�E,л~L��UBM>���@�N�c�#����7N:�$F,�r�(EeqX.�D׽��2q��H�#�J���2��Fn0w@��%o���WDȲ���>��֧m����f����H(Σ�n�.�	����-kǢLP'ʑ`���x�(;Yl���+jf��I[.50�-T��V��IZ�z|ښ�7n�hKze�J|9m��������*��e�J�6ƴ\N�(�}�c�G�a�}3,��y|��c��A��������d}�������ݸd�����BEB�8��s�z�42�`x�Tr��Q������>'84D�W�a�ߣ��4�:�J��������i�g��rw�U��b�}���w?�<]��XQw��x344�0�99ǅ1����ii~&�{ ���7�ǿz����Q�@����(ڇ���l���V���g��%	�`\հ{֍ĭsO�Łs�UM}��Yn<�y��r7ѫ�����:���_�� ���]!k�c�+ Q�����t�O�}�	����0-�t�Z`�� �Z�	�hu\|�cE>t⍳Hy�j��*B?�'`J��J*����`r5-4t�k��h�_��z#�f�=~�ok���g���4� \��ۯ�j�rP ͜?�%P͆���Z��V�a#�L 2�G�dϯ���g�v��l��w����Y��¢^:�x��EN���$�`�;���W��~���D,���������ܬ��$7���m�;��x�D�" <�ن��g�_\;�����O�ԙ�>_}v�S�G��!��Z�'��bt=`a���]CS�.K�Q���l��S��O����4���]髰��Q׀�JX�3ss&�w9���f��� ���#/��7���;&�(��/�ݱ��C��IB��n�d�g��DJ�|�;��n^�/��J*}�kV_'(�Y�n+����zQ�P]�6bPҞ�~^��m�S�m𘃫�Ù�-�j'2-/ꆆ�͸���HM凧8
b�lz�Ns?�ٌ�_�4�<3xV�4o�n	�+������-l�����$�J�6�O�~a����<xR7aX�R?�:�9�S֤�`ܫ+�ΜԄ�RP	o��1����X?��23�:��$$9�N5��߬�+�E빂��'S/�O9 �p#��������Pwwقn/oq�л�;sq?�i��qk����	�
��X�����e���9y;�(� R՜��x��s=D�o���$%��Aʹ�E�p����&�=�C��Č�p&�,�JM '+i\_��
_� �FE�]Qs�ٻZ�Qk�Ў��X�`H�����Uo}���A�5X��R��g�%� �[
5����; f�id��TD��z$d�g��A��c9�9jj����3R&rZX�� ]�=��Uwb�׌]{�~�b�^��B�\M�y���6����źT�9�d��_�wH.�\\���,��T[�d��U:Q�ݖs��'&p/TD����G<�NA�gX5lL�'��vW*�]�t�y� ��ٺ��xJ����gcJ_��Z�_ӛ�Os5:����l����W�9(�C��z֕�_
B�L7s�����;L��L�6 �3s^�8<F	D�t����]�Wӟ$�����(]�7<�Р�8*�y~���sU=w�;�?�ntp�M0�� ��B�|��_�(��R� �1
~@���~>�y@�"�7���>+EP�;��|�jF�G��s�]}�����M��_#�yk��B%c��e�)�҇���&v~��;tz����߀����.e&���ٯ��_w[�V�ヷYT�#��"�}�J�����:�D�]W��X��r���Wx (�aD�À�9��/��>O����X�9�g��߳����+��V�uw�qҺ���U�yE�l0@pc����=M�c��>X��f��w6�j���K�C�c[J쾜���A�j~�1.�LEЂ�)[�~��.�ͯ�/��D�q7Y��%�%�����FZ&o3~�v �&�P���j����D%X�N�s.i�?�B����փ���s&sBv��h7(�l!��d9r+��E���Q��kc��S��n��ΆW2,�&P.���i�(���QtH��R�P숞!T�d�Q�_��I�ۂ�T?te-����V���m���&厮�pz��P=�t�=���8�[�#ԧ���=�J3,�8�V�ْ7!Fkp��Q5jw�U�P�Ի�"��D�r�����(C_�M2���]�m	%��\8����l���3R�}B>\����R�a)�0��MVG9#��j [��#�/��:��?��^l�O�����q��Kq�@��V_>o+�_�[dr,�:��b�\��{�9�W��V��{�� ś���z���<9{����@x���ǋ�z�<��c��0+�7U0��-t~��M`כ!L��Zg5�C�[FErK��Ѱ�������&L���#9��N�h�o�_{��^(��|7x���]�Yw�
_�>;g��V7��Ǩ���g�I�E*��6~(�Q��w��r�Fg⼤���N�!�d���Q���N�5nc��E��SŽ���4�!�j�:�nYC
�b[�}�z<�ҖX  ��+.7@��1�{kheXP�o_[j�AH�&�j�y��V���Z^�� �SN�߈�؛�,v��w�)P8O����� ���ᓚ翗.���9��8�UL2�g��datSԺiD���
᮵���j�rӿ���P4�w.t���{�%ֱ_,�~#(5ۉRI����Ա6�?X�7�V2yLČ�fϋ��_/�b�a�[����l��5=$r_a�2w��;_hp�c��i�k�I�������yaXm^t0WEI��k��B���ݬu��e0�G�8DC� ?ARe#}?����,�UZM���i�U�tW�2R��v��jQ��Ai�ݟ�VN���	_����Kf��8Cs�,e�sY�� ZQ��_�6/��d����+A^�sӋK %
,�r�@��DC�����P��~��4�3>��[�Ĕ"�G���{��ū?W�f��4;I�Q�nLdCV�I0WV��Ua'k����ռ)�Z�:�f�j�S�{$?�y�!`����}:8ٕ�r�+�1n�a �������@i_e#����i_��1,��t�o���$��� �R��?�%Fp��R}�:�CY��Ք _^+�Τ�'��^�UyB���!��,���3G*<��7���N��>��aeUР�>6<a�Qo{)bf�-5���0+�8r:�����Ĕ#	h���j�m��o��Ù���V;\�x�#I���C�A�O��24"�x$�Z�����Eb���q@�v_$��BB����D�B�°��$wr�|+��hn5����bx?t����Bvp�ѕ��,����;��M�w�<��`�
��L°F��*q'È�� �*$HK�l��J������=Qd���W���ܫ�Z;�Q=�Yr�Oc��
�I+H�����&�a2�����H�Y��M��ա"#�-S1��tz\��1� �\^Hr�� �5A�w>=N:�w��I�4(�$:@N�}����jT|�p�G� ��	�G	�5�G�m�N?XmBz�Jj|��'��|c������ 3�`���K��;صؾs��?w�����O��=w�`I������p_��I{(���א�����n3?��td������k�c�vr��ؐ\��
}�Ĳ�����\8�5
w����Gs�\+�xu����Y쓹��Q�vi�.��1��ĭ�")ATj!_�Ɓ��ِ���՞�1�=!t���1&7��3z`�p���r�n��t�����TaC��o ��-�mhR2�\��nk�,\�%��䋨�r�t+R����F�`�6"�L�u!�
^��{�(��d4���U�G�e�>��q"�w`ô#��ܖ��Y4��qK��p򍽆ho��~ �fݹ�����3Z�b���hy�G��a	��a`ips˸:�T�d	l�]�F����)���'�t�|�c-{3�ٽ��C�3;�>,���4�r�����*q�<ӯ���#��6r87����a�����.- � v��㋋���3�]���J#�)�@����|����/q�7�J�����[6m�!�w(��敻\��GC���k��z8_h%�l��!�4���s�5.�_����<@T~�)�R@��6J�\.HL��6�J^=���]�
|���j9������'	�E�G�#݉��m P�+I� �BR3^.+�O3����T�8qFw��V����	�B�m�-V��P��FpwbZ�v��+5}���k>������_�8��6���a�|�o�(0_[�2�P�~䩶���w��ža�Ќ����K�j����:�Έ�'sZ}������^���=�Tz��w�<��D��DIT���h�Y�e��+�|l0�^�*p6����2�%���E<�XM�o�[!�L�E��X��rO�l��r�m�3%���<{�қ��0M���&�x+�uqG��>���&k�fSuj�8�2���3�IY��TX�B�%-�sd�7�:�_^�����$ ֹ��(G�ڱy�3t�A�1�WD�qʐѶ?�`��cƓ�	/�pf�/�v��,v��	�A-M���ͪ1��b�Q��i^x���u���{��I �Ƕh�j�u�ɽ-�v�؉��-���(sz~�UeǍ'���/O�M�.�?��>�j�]�Y�4��*���pOߵZ ���v�����ͥf�e�	ʔO2}]��`Z���C%6�й4�O�F˿�^T��81<U�L��0�]���"�U�QO[,1F���7��L�¨�$M�\�殒.��(�Ui��u
�.���m1�Г=���ׅ����1'ix�ǿJ�f�e�zWU()��:J:	��8�X��v�;�U�=o�Ha�k��:������ٌpOZ��Z!�����*5�9��O��������:j	%ZѨ��b�K�*ݻW��2��\�P~6�ǈ��J		���f�c�m�˘�^�c x��7�^�Vbi's�*+���W���ֱJ=������,�ğbG���	�B�`k'Q��ף-�h�1΁��C_�5�������k�6ނ�� oCȄ`�0�*�%�*���@�:����+{ ��A����ry* ��D�٠6'�5wm-�����Iys�ۿ��B��+��r��%c=f��e��R`�S�H'�&oo&�R��JL� �4�	���7�����@�UP�@�CvC�`�Ml�:?�'��� �F&XXV {�cTI�&XRpo/+��Y��j��>�;e��_\��5��d����L�7�^��@"�c�,">���j҃xZ������ϻvHB�;���#��/�f�����9�$���#h�����+x��O�ImQ���qz�<���dmB(K�]�nc"���6o_a�Y�|p~���b����eTI%J7���
7��~��i��k�Ѳ<��G�ˍ�"����D/t�fl�pd�ђ�d}���^&�;���|�V�
��G>�X��i�+��3��^c#_��zҼ�#����"9}�(i���p܅X��d�eB�1��h@|�s�S�W��+����Q�ځ��!UY��5��ə3f��n��x��,�-���ݒ��e���c�h3������ЂƮ����; ���b !j�1$+�+ �v�e�z�%m0���̗Y�25taںyB�j9'�#���9����62���m�vr�\p4%� ?`5}�M�h�7�hY58���8�B���r��y�<�F�zը�U�3��p}�.T4o��7�5N97�pt|w5E:Eq���d��]M�i���=�GXMRfbYT-a]��<0���J ��ա��?��
3e%���]��S*�W&t�T|\蘂:4p 5�o�!+��(�������	�P��M��Ҍ�b���\t��FB�ш�9`��En�lQ�8J�a:��X�Z&뇗�*&�9h|H�DÎ���^��#H��R�4�Y1�b8��I��S�<����f�k��5�{�q�$PE&Z����?`;���^S��]�FL3+.�1�Uz��6:� {����\��D+�]�-_׶S�OFfO)��F�^iɻ�x_c��52���d��4�\�����`>Aݑ��f�`&�c���0��+���Ǖ%�YʞZZD��O<Ƿ��_h��|����Vf�H�NX�v�dX(Y�,xx8�n�"\�����刭W��8��~����������� ��I��h��j�� ���vS�_������?��e����Z\���iE�n�!���/�ܭz�?��zטNș�D����W���A�cD�/ݸ3&v'�d�������G=�ѐ��o�΢_�G1�5��wpx�S�	=�-ՙ����<Ƃ]%#LwBx���RK�0�����i��q����&/AwE.�����2ȽѤ	��ݛ�����X�������R.��-FӲ�bBb|#+�@)2�0��1����*,֘�Ղ-�] ކ݇,�
��v�k�9̦2��%��uw?�����@OT��x�B�k��� �4�> Y��신]�A�}.������;��~d���st��ɾ����tȌ�`��'���Y���G��7I8:��-7�s]��i�aK$
���'�2���)�k��P`���Q4�5ꨂ�Q������]7���B��Տ����i�~��^U~�S��H��^��^�+�/$�c8-�.���C\��~���.-r�<0{�ϥ��x��^���nF%ѳ��t_�u��Y���\kml2)�7���ͻ=�旨y�E��6�ۃ����	Zл����@�uc��K�5?+��ߑ�OY��kS|Or��h0�]'���'��s�SJ�#}}�g)��ܦ��jB�S��=W�ӹ������٦��Xl>���(/8�0�� �q!Km%"��OǼB4;�o��˧p��
U�$J� ���`�y!�kjy�]<&����VsNh�VM<���H�e�o�������dE�8���x�#n0 �Vw�S�˖?�ma�!7���%��S���O6+����\.6*1�/���yU�ڶ�q���O����N� �#i�)���Vx����P��I$2N�t�����7_�W��A�|s���0�x��
e���8p��!%� �1��j���gQ=������P��V����
�fSɩ?�;�А����$�B���,�Fҙh6yw�.:1�ʇ�.�-�,�<]�OW����g��]sAqf��hO�M�!�%�?,�v"P��Ҵ�O��V�.�HAU�5-��� �������c!G�����X�敩�fV�֣e(-��]6�Hbjy�������C�.�Cu�k
6����_t�/.�Ya�<����� +xY�F�Ug/���"~��ʘ~���H@��c�bc��1���H��++�Szo(pI��,�GE������#�jksJ.ӿ�>EZ>��s�j�날�ޒ���5<�^GW��z��D�f�Ω���������^j"߷9��s��8�ވ2�͂�Z�
�V� <�����h������Ys.'�m|P�1��]-�~� �����Ox<G� ��&G��z�p�L֟�T����Ώ�!X��Ĝ�
���M/�sD;N�C��P#�z\4�f)�����0��$S��?���/ I��U/`~le�j��sR�Lz
�|.��<����v�~��pĊ�e�˞��ຜpQM�^�%��(���d����ƫ�ɤ5��[-�h��E���O���p9���ð���U��p�?����ŇF���)�^�*�4li�͋��N|.���'̷pz���yd~��w�U&4=H��`�Q�C���;��-2J[R�)*摱D3��r�l���"�[��Pֈ 0�q�Ha|��
�Y>�y�rJ�w�g�wDĞ��P2HY,yۺ�>MQ@�[���Qr%�8����T�H�(s:H��e�����(�@��W�rJ|���85\_���֟� ���|�T4
��Q�|��9��s��N��u�y�	pû#c69����F"&�	J�Y�Gz�����"�Nw��m'���4�xe[��鯡.��b��O=#*d$}ߺ2Q]M�^"�tl|�T@��WsoZ�`!D��&h�\�M�����靽��(+�"�D#�lɍ�{�8��&�6�h�ag��z�s3�9T!UPN�]��N;i�;�*b"��J��^�$?	<A�h��t��q_�C��r�h�	a-��C=J���7�%#I���r��:d�u�Wy�j"~�8/�/ zW�и*�l�f�� DJ0����ж����+�>)�^�oQcz�.�Bǟ�j��M|۬ҧ�ێ��1��6��зm'���5j�2�X@���^&��ƣ�2@�}i��"2ܐQo	�R`���h��Z��R�_Z�Xke�� ׳4'�a���Ča�VM�� �|����3\�`�U���=�����.�K]�E�q���A��j�����׀����i��K���)S�6"������&���"�^1�Ԯ���1�z%N��y�{�-c��`��Z��������V*��C��n�bN�B�����q�|�� ��|S�X�V0��SY�d�e�P�4AC@�Y,�a1�Z<݋:P���/��Av3OA�?��0��̂�9e��%�!�B	nl�\�y���fe�B�j��f�1@ǷyW��d���a��������w�����M���#�c�(7��*�	�$�7�:u=�p~؃�b��6�f-{�mܩ���LU�V"!�6B�K�u�suΔ��IJ��[ ?���c��AÔ~�T��*S�QJ9��ATp�Kn�X���;�Wc0�V�ې!�*`��W�y�#z ��g9]e����u%kb�=����;���RW"RP3V=�/�1�sK�6jn���z^8�R���ΊXa���b_������� �|�{����d����B��;�X���Dq#��!F6?�ͦq-�B8�̘Z�8��\��K=��6���n�~����hK��[������4��b�Ds�K�������f��H��B�#���+cx�u�#|����>�xy.$gǸ���a�C�M��f$ɿ\�s�
���>��A�r���X�#�z���4�$������M�@�-B�sPq���Y�����P��YZM/���ѾQu�M�vc�W@|�j�����!>�볭�t)��~��{�t�f��[Y��^>�*����>�8t-HM��l���D��odb�p�H���fZ���F��D���wT��5���*"8�a;������yw�6/�%b;��ɺL��8�O`��/��%A���VC��i���js�*
O��뭇Uo�jK]ŝ�n!)�7��_U|�l-:
*U�S^?�P���+��� ��G(nO�;�~�xGJcZ�b/��̱;�pQ�όpHv�,�>b��� �_�>���8�vL���J��RX g���ފ�a�j��3�:'�e�M�@_��O,����wn���J�G�S�<����L��L/H�˴JY(��	t�^�0�]�}��uv9.{H�d���2b"�����'
�?Ĥ��-��:�W�K��0��p�]u)��J�� ��qN�y��E�(�XFw�6H�ˊW�C
��Ǭ�9An�~1a��N�5P`�������9�b"|n���=&4.b��!����^E���N�y���������+D�l�J�X77�ي>M�i\U�xM�Bb
Ѳ֐ި����j�,%§Q$E�I��'�X�98�篗΁ Y���b4<��E����%�ޓ�h��,3L���g�k`�ў��oD��3RK�?=�1��`L�M�ٳ��>e��=�'��֨�D��8��Unj��]8�{�b��R����o4��q�Иs�(�I��M������Jz�T��go=lL�jK��"m`�Ug�޹u����x+����O���S��8�~5���A���O���
�����p1���b�x��Kp4^2�UF�Hi0L�)�D�	E�xV���eI��xZ�%K�"�iQ��4ѫ���mݖQ>a�_=���>��fĂ��U Y�~[��z��9�����r�v���tOz�=Ux?��
�R�ٹ��q|�A���ad�f(eF�S&2*�b1���P�Ԑ��}���ԫQj(�2����N*��"D�Z��5R]�?���	�Mk�ʑ�� ?�1�\��j,�B܀(��,�>*��S��~�x~D��G�,�+t�u�0e
�}�Yг9a�^c�9��li�����G��|�\bB�rɻ��$`Mb� �CGy��U�U3�sK4:� b�*X�X���ݴ(%je2sL
���[�5�m*Y���4�ji����Md�"����t���q@i��o;˭����%GR15��T�V��<�W'J���r���P)�����UPs�����m�>���t^�$s�v��\+d�K�RDh���v�.db�Ѽ��[%.X�o�
�>�x���r4���j��������K2o,vb�>�״��)ׁ�Ԥ,�~���h��&����w�[r�0�&��
�m5����'&UwG!����"�+�b:�Y�����[ġ�w��֡�bo8
����&����Mja�l��3p��hX�޽m��=ƘJ�P[Q��x�>����(^ax|)z�P79q.��#i?�Y��������,�Ћ�UoH����Bɧ���{^�+�)Bù�*
�������rmY0�2���3���j�a��
�X��U��gM`�F<j@�9-:�EN2�!s�:�,��b��1Θ�i�UP}=�ڼĲ:C�n~ǿbYז�m�C�I�nO��|��F��2iw�i�� ��X��T��7���ޕj�'}f��fe��k��>+$����ӵ���"Jc�3��&fw:|����sE����� {�W�S=k���q�H O_����O��kd�ZK/�M���8��������0���������G����$�� �¼
��=fU`��!0oj%���)�ꑦ�vQ��k��YD��9�����`��v��ŠNM"�k��+�"ݔk5���N��Ά��>�0[4��RlS�I7T9٭���QS���ʁ��"̅=ؤ7��2�(�
�^�s�NdqOߨ�}vT�����=(w�y�@=���yk¾�����LZ��uZ�w0�7�|�����ލ�X��������*:=���!e��L�}��������>�Gc�[Y��n�Y�U�ÎA�!�i�c��H.<��B\jū��¶��lB<ѵ����#-�d�r�2��u�	RP�6�N_��A�9�e�#�呢,4'W�{�E� �ww�(l�V�B %�Sw� 8���t��H�`s%���t���ٰl��Σ_ػ�`���7	ļJf�ԉ��mJᮋx�,;h�����tl��~Hiu��IGF���E�G���n� �}~��|oHMw}g���5;%���H�R�ٵ�i 	��m3���JEqW�!�87i����c�p��nM�K�m�y?~	�:���j{�@�nGn�P�}L�����ވ"�+�r��>���x'���$�k�A!��;�'�:�:1~��u[�w7e� >-�p��"S-6a�F����� ������=>-s�[гd�$4�I�� a+�Q&	 ���+}�`U�d�QC��ќ>�_؃�[Ո(��C5��>M$��0�Y���zY�����̨�	��G��[αuGW�v��J�ot�/"h��i�]�p�jc����$��by4��k�\�$�;|�Y�>���#q�i��ɧT��iD� >v���J�9.�(x�K@/W�f�zm�vm0噽#�ٙG�'�Ky�)����LV����C=�6b=♵@F�'�ԍ��F��hi<�J�}��%��N��S�b;�.b��M��ZR�fMI������SPl4t�&@��IY4O�ŋ~�r�~1�UĤ[�e6��}:D5R �.7]�{��P�㎔b�5��[���PCWZ=7�q����@��1����S���u�wKQh]�K����,��5����UQ��Q7��)�)�^��W��F�^����#�޸�Rz͌�x>�7��ܥ�S4����wbc!v{?-�0jd��b�$YwFOZ��e�������GU��y�I�M$N0�\/*�Eʳ4&��k��&�z��a�N?��#�� ����'��>G`.+r?�o���P�a�̻�4T���Ua�E �P�5(����2��Iՙ���dJZ�O��>�	S+p:Hm�R�l�l)T�D��)�}A�#�{X<x�l���b��ò�1�kLBF���ǉ��OSż�v��
* ��`�^��csacy;N�z�Bq�ڥ?*��������0f����d���K[Y��W����r�K�*�L�W�z���DL���;L�K5��8v��
\Bm�uJ�W��}�/��S��#YSt�9q&F�x�Ɏ&��:@��L2�S[�	F�nK���9R�e�x�S��;��&p^�4�§N|ߔ
�����&�F������X���S��G�"�׻̕����+�B��'1�&G�F�R��
[>����{M3X�����v�/�=�8��#2�1�)3�=�?[�WP�è��ڜѰ�l����J���>��'>	*�9J��	��3�������d▞Ku+kB|ǣ'�H�E皓�.^s�$zm!��Ěb�E[��%{�e�X��"�NO�0��j�O�i �-`�-��]�?c!'ݏj�K�֟�F���;5_6bs	E�9�(��!���u[���1��[�N�Lj?��lE�@#�?�D�Cj�"@QO�/5no[\�QYs�`��A�@b2+!�9I�Ѷ����]�?G}������u{��g��W��w"L��Ġ��*�0�� ����a��R�U�@E�P�fk�*r���K��v�H�
>�!���-m>��Q�s��>k)�-~7$^�a�U)�H�\L:S��e��R��[�][�U�w�	D�\�kB�ք�%"N!Ƨ���Z�x#�$��z�w�V���a���B@��w,��}�Y���L�W�s}0�B'��i	X$�I�)���Zfϥ�����Z�M�g�R�f-Q��]4�����)����%���{w��U��x>�vf1�I���>�N�z�>Zojb�d��,���h�Ϟ~�)X������մj�`���&Z��Q�ooC���=�uZ6B�?�55S6*�E-��EȚuq:����,zψ�6<��d+t�n_:,7��~��wPJ8yI!��B Q�I�aɎ`�r�����	m~m�XU���5+I�~r�z�IŇ����kVl�����I\��Zm�Kj>d"���<�q���S��&Յ��&"E�	��y\���L����d3�ݍ�r�Niz�w;H��$��fH�{��`H���¾�)���kW������L-�^�`��L�A�A�#�3���ayX�1�}i4d��t���&���n�8jإ/�'EjB��2]��P�ە�fW��# F�.pd�����Jz2R���Th���f�_l��қ$	J������"�2b#gU|��[��-��[��i�D�Io&�u���y�J������z+���%�;�O������)��	���@�*J��$- L�9�)���hg�t"n"5쐞��T{*�t���k���y�n<���m��\)=��&)��+�P�}�X|&� `���ݔ��̔
AE$qh\f�s�#Ng>�^T_��vj�=nY��7�����o6�;���m����9W8��~�S����Y�<�!�-���W~�Fi�[�o#�t�{X������6c�Cs�*�؂�b)�P��I���1�)�+�E@�a���!��&>w���nd�)}R�>7k���o[᾿��?�EI�bw��FyÉ�fEa9�+bn�	�����e�[�+8��H�si��$�z��"������:�����,w���ea��t�!�n��"�(�P�8(�]�I�-���)�Dś��'�	��ߴtK��qW��E\�V��=�&Z�+/X���^|D������p��7��V�� j�v�~�bl,��\��}�jY����ӳ|	��Y�pg ��rqZJd�� $W�*�̩n���	w��4&4-.�=��1C�b�Z���!���������ѱ�b<��%f��x�6?��u�ut�lÈ��Y'�$+�w:b�������3���n��oO��%zp�NVKyZ�$T[��"���+\�u[,�HGGߤhA��/�mN�?X���'N͸Q�5�K�l He�� M��� p�������D����tn/��sXcِ��0�\rF�aEtA2�3Ѽy�|q��LI2mz���wdO�+� >~�|tJ�ˡmG����4"��p~�Gj�}"��`m�q���O�r���L�Ji��#�,~�=0�*�9�'d�m*��$)V�j<_~ ���i!S��g���S� g˺�ۜ�?���q��,5P�=��G�.` ��V�������]�=��p�A�*�\+�r	�����RDl�J����y�5Q���}���'�w�����W�@z:�-۩d�w ���C��v��u��	�H���xT�$ݗ?ѷ�%F��s��]̘���q�$�N�3tn��)��h��0��
����S
��S�2i��W)�5paJ��Pgc§~M�g���H?R�հ@�N+ğ_�{�R����Vu�:�z�m	\2&�3���I]��]X����Gi�W\c��͟P(��x�X��t1RBR���aʄi6���Z�; qa�����{}�|�Eh��.�s��U^��³3���Ǣ2�z���=|[l��~D�;�z�<���Qëv O5,�����a8'R)e�c�_ڔ')���
��E�FR⒄�r�(͖O��uW,ء�+O)�
�R7C�ry����}�턭H ��#�M�UR�_��쒩�T�H�_~�B���j��H�J��@���|뱱;!;����r��o?����s,�"8YbW]l�=wU;���f=�J�]�?ڋX��p�L�	�414�`��;�|�'vF�͵/~&��0�(�Df_c����7�,�_8�Ρub�.�X:�4��Zf1]�?�F�꠩
0�W_ac"�q�h]r%,T��A0䒑�����G��p�("� �*bN���{�$����Φ���
V�����^9�v�	CMaP�4�a���3�d�y/*�������n���}���t�fUJ̫~�xcA��2Rn-���.�Q���U$)��4�|�R�@����N���g�J^쥧�����ٸ�a���F<c����U��ᬆ2d)�g�����%K��	o��f����ƍ�����a�sS�_���R@d��2,�q�Z�����`�'���%�/:�5<zϵ���*���ʷ���Zp��
���L�5������F���%�>Yv��0�k��rZ��߫#1�ͥF�Z򾡵�U�����#�����Ǉr}��|}�h����*���F���P�*((�(��*Ӹ����\aR�P�~��}����N5�����^�HU���!B�i{N�T����x�E�>�j��_�Ev ��&L���t�DJ�;�4����*l~]����o�BS��8�{_����Z��H�2�ԠY�����[��]�9Z������oJ�%ȧrh��ݔ��!��̖�(lU�z����&fl��mFܮ�ȄiЋ����d�,e[�#V9�R�tL�͞��7ƖS��}rV���Ǜd%'p����h�g����u�ܘ�焊S���5"�C����~�_ׄ�)��.�6&����T�2���%�Ԋ/C��kH {*bK��)�?#x�7��M?+��b:0�]�r7�>$u�ɏ���m�E�����`��r��kj��z��S����B��haze
��ֽ����]M������Y��ҿV�N�T���Q�;84��䇢��z��V0R������{mU���(�vұ�]{�Z� �<*Z�r�>}0<Kqb���*u���`��u��fzOɾ/����ul�}\/��K��%��*N/^�D6���{�]٧H���?6��L����Bj��*p�(py��t��+��P��)�{m���	���� m���l���_����&����vTnz�<�
��eF�5g>ȥ���������X|�����f��0?�F�����K��I��;u��?���" ����Z�	؊ ,{��N�3F�o�%h�C��-X=��<�k=q�9P�O4�̈N���[$=q�����������
�蒧$�Gd�OKۤJ�eL����u?8l�2z�֔�,vD��F��鐛�(��g؎� Շ�G&��#I�Y��	&RO�Ʉ�Ϻ^��ö���:��/��/*��i��N���w�ܰؿ*7�:,�7v
9��f�KU�뉟OBz�@�����C��_V�����L �\	�����5B ��ͪ�˔��)�CE|֎���hvvy2z_H^8p��Y��Ş΢��SK��Ό���|���/����C�>�a~�;��\�!���j�� �QY�Sh\̡D��;
:�
�����˿�?|2���.TޅGp��ȱ�p"3t�Y>�Ip���hF��5��׉�ń��<���]�Lт��mD�W]�����`����!�f���횾aV�%�
O6>����&c_����V�Z�����X���FGu������:G@~��\\0��/��Ŏ54�L6�8������0��JR�"��z��7��sP]�p�W��%��eBր�)����6n�l�aB����nCI�H�?o�h��?�]��q�r膼IR�扒H�w������we:rT���3t�"j;��&�t)��;�=�K�+�{d�b��I�XlҬgo��2����1������ƅ@cI�⏻~�����d�8h1��Qq�3}b^+}�ǽ�$ 6���Ƣ��+4Z�t{H�gU����a��8��'M�C�������ƶ��̰f��g�>3��K#I��SK�V�w
�[�ڸ��M��+[�\���5����U�����<����_P,�鄛�Ͳ��B�}�t� �!��7�^2Ѝe�>�s�0�FN<�&��$Q����G��I;C��<���IS=��C s��Wy��چ�}%%1�T�S���Lv�`u��l��a�^P�Rh�}�A��������I)
��i~�9n��#���v���r<'��G)���m�R�� �Q,�FS�fه�bÂ8��Y�Y��Y�څ�� -8��� ł��o|Dh9|��-��Uڂ�S�M$
�XW����i��A2��t�l-
��-r�A�����
��9$b��uc��4���S�}H Z��?�:L��� d���8E�א�޳��0�H\kU�}	��#�W�g�UF?�#>~��}R�\����c(i���<��{7���i�ɩO�RM��S]�J����*�����S�����/g�7�̣|c�	�����0N�P}»U��%vd����u%2�[?�ف�.tݓ�{�޾��U��4��/��/���di����}c��7\�r��e�
p���׏e?����[&7Gz����o� ��HP�I/O���@O�s9U.T%�i����5	�����3?�z����䊲t,1�ӓ����#�7ݚ�5��:w-̮8
�q�:����>ޔ��a��@_�\Y�=�J>(g���^e��?�î��*ǴVm�>�ʽ.������,�})������_��iPd���τ�`����}�Lj���]�'9 /G�d�0�	 \{'0��*�qj���@�P�-a��T��W�쭽��vg�u�q<��*�*�M�6�0BÀ-P��Kŏ5�
���V�Q�o�!Ѽ�r��q��g?:r���~�e�dC�Gׁ���`w�Y����]��u����4��{������AnB����u�2U�"`zp�j�W�6I�.�T�x��0��~W=��c���w�	O��\6�_���y�{�yR�6T�IDl���	yѠ67{p�'�L�������煘M��'O8���ѠqN�j��:���I���a|'@!��ce����jB��b4_��@q!�Fl���q��z�����$BfX1$�*���53Uf����/P����ʀ�H ���ޑ�N�q\��-��9B?B��ڐ��F�������ڷ@6�yo>��+�DhKz�����+��?Xi�.i�|3� >�u�WQ��o�ΖK�/�Yc��3�lX�b��E��,x��x8�:�߹w����7#w^$�gmW��bO�љ*k�A�W���)�G���[7�@�x5�􋳵1�[�"�����[p�ޙɶe����f�,�~ZROd�cc�U�z���ʥ����C��ѡ�4R�����Y�}�3H��ݚC5|��/�-r07��?��1}	_-Y�q�UI�M�c���8��6��1ڳ糿Z�֖��m�GV�z���g�+,d�X6�Ƒx�'�ͼF��_��_�96��2q��y��/�M�x��D)�D��a�,1�|�R�z�J���1�u=At~c�'2��X.f�^A���y.pD���fnN�� �(B]x|���$��9`W��Va��vC�W���7���)s�{j)yU]H��1US��PP�m�L�`�<���k4��r�ub�Z՚1��X�A^rNf�_4����m�6R,�Ow,��*�U�-� H1�����M:��o0NT�2��z˚�E%ᑒQ�hO�W�B��Xb��M���s� ���/�w�q�����+���/��% "�㸾��Q[���S�S���~�AX�D� E�哦��	xе�Y�f��9��MA����ׁIV�d%�0�6.�Xi��8�H���[2k�Q�A&�������L�8g��嚱��bQ9�����ӭ!=K�q�V\���xU�ʎ���� �h�ɪ��by �="��2"�C���No�|GųfS����#4�-��Y,3y�˔�y�h�6J����	�ʚ��.]	rr� ��ۏ�aU��]#�ؘ�D\�F���Ӻ%?M��y�QD����9�`��@g ^��'�D���>n��\Tm��L�i�����݉ll���r�g����6T