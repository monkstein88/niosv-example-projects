��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2���f�[��3��}(�^P��$�3�ۘ��%��A�Qx��C�EQ@�{�y��-	D������[�TL�Q��C6�74��7j���p�#�lM��ާ��3�k��!�
���n߳����h/Y��G_��w��"4�0���R�W UW��Q�j�:UAYQg�e��m}�$��s������Sڷ����G��y��Q!z�Eh�hHW��e̓x�����Y�)�>1�I)���᫉��æl,7j��������M帻_R�)g���M2N��K��]:��?��YZg�!�)�p�`�3<2��xY����K?������3���/v���6D�t|T�Њ����r�OUj����:�pQt쁭�܀���>WP�:%K��Ӱ@E�N��9s�1�&4��	7�j���}�}��\x�QD�f(�u�ۘ������T��>/�7_��g��/X����:�|��mQʃ7t�h��ޢ��gJ��71P���`��[�R_-��z�i�R'���/�w��-aT@�+
�e��y�Dh�	$;��I�k�G���{�u.�c�����\����|T,�!�"*H}x��ק7v�[F����=����?]\�P��Myֺ QS�8eG8Mm�m�Q���pA[���)���텡,��[���ߣ�4�Q�LwМ؝�;�	�!@\Ȁ�߻�����y%�M�����K��3�e9��C��t-`7U� ��	�NFӿ��`M�����]���N������𢡊��]ϸ�s�LS�����	-,<gܑg�}�aH��~�{��V}�Hv: 98î�3!�*ߺgV�w˓�6���k�D!��@�a�n��
Ё����}-×~E}���y�H�;`{>�G<t���$���@Y\�`T�,�W4��K�W3�d�Fi�Y��ּ�����Չ�
��V��_pߢ�u8�j:�=%��-�H�	������Tߘ '�IP;���aPY���5*S'��Z�Ej���䌬�Z���_�n��f����)�&nP)�i�L���R�<�֧
"֞�&7Fv)u��z7ҟ�la�ET#'�Bv��x�(���Lu�����>f����=	թIV*���A
T��.[>.}1���S.����@��K7Z��9d�^���
�.?ɘ���W��������, �3�Fn�Z�y+9[T��x�� �Ǘ��1���3e&�`ވ]�s(��TQ�����&*ᣇ�[!y𩚛0l���ʭ}PLң	�oM����;A^��̀�J�9_�z&x�-g3��Wϋ��PQG�f��~鹰J7����q7%�ҟ�'2K&��N����(;�"E��ڭ���gCrx��B��/��؅!�Dy8wMZd���!�������>�|C&����2���@ ����U�g�$��<�5��]*S��G���Fb���,L:��[��_GT'"�{Ԥ9ml;��n�&ϒ[���$� �r����٭a�o-���2M���ee'������'�]Δ��`Y/����W��5� ��[:h<g�v��#��Pܜ�H��lS/�#7������Ж0����޶��1x��0bi
�`����Z;)�b�B�n�����fCh1_&�l뤂�rq�6�۔��Ai	�]QK�VEɏO�G�q��a$(��nm&3��$�I���D+P�;��� 9!&�+�ɛ��=�����C\�R���d<��^�^��A� �0�4
1%� ���<���b[%�#�ʉ��X�|�i�J��UK��H���{r)����$��J�pD�X��0��^�=�Ek\�{0?�6hï�@fa@�˩�=����ʩ�����be'c���x����+�ٶ�{Z�3�����x�F,7��}�(���Sw���_�e�1�6߈g� �o�~A�A+"�\s�v{E�oO/�#����{��$AY��@Cԉ[��Z�C|2Sw���aO�7M��+��>ȼ�s�jNN�оZ6�9��w	�ւ��%$�[�\�_�I�%4O#O���<��<II5�Bc�����\��c�}�,BX������S��/Le`Q���ҫ�!-��M�'��!E��L��'~�$w���i�_�"<	��t�D>�ٙ����d+�DyAىr��/-�`;��m���g����/~��k����|7��d��p�"cm~ע�"�~�M�8�k�����Ď�?�?t��+�W���L%��Ҷ�0���Q�i!<�dy���A���0���PA<U��0�����6��^i&Ɖ#KO�Vq�����UU���s�:c~0�Ul\V�e7���A��AN�����d��V(J��D��"�KMC���!S�a�%�������d:�ON�
�$#�d$���(�����I�4��nX#�=�s��\�7�L�P{�,��J�ے�[����H�Y}�zZ�X|h7����`�c��K6>��ySthY��e �j�-Q?�0�L�m)������n�_̄Ȳ-���5�eS���m�H��4Z��t*ɰ ��ݪO�"Eu�f~��K��"������ߗ���n�ș�Yir� �o+Ca;���UV�p��wQ�"�y�.�Ս�B�IQ
�*��\�������ꌼS�G��?�!�p{���+�ի4�Fo��x�%�1��u�JP��./��]��F�Q_-єT�.1r�t�S3ڱMp�d��V5�f᩿�F��>��0�1?ei7"M�t�K��^=x�(�����}�C:���B�z~2����NW%�3%�F�֏��٦�:���=rꉖ��o.��a_���ӛ�1�@G6�8%A>�?��Ts F�/�&}�?A��P��֦����z�I�O:�Y#�l��*�y���P��QV2���1"���~�اHb��S��Zxx�I�NC���ƴb	,��u@v�&�0Ar�۞ɝ�=��xϹ��<2��|�k���;���K�[x�����c{�Dz8�/��^J���`�iKw_/u �x8 ������<rн��> ֗_緌�C쬣����bh��R|�9��_��҉�����>���(i�I	�_��4�h��&�0�0�[5��W%�쯷Hu(�
!Z&6�j�"A�!��}�\�tN�����\����0&�\��I��"UTf+��9]x�/*dJdR�O�fSC�����5�����!��׷t�&2}���bK�0�N��6�OG�@��
Xl�O����so�� �Kֻ���v'\Q��A�Y��V�]��	��pD_y�ĵ�x��(�(�%��w�T�`��D3��W���Q+��z��6*��k��1���o(j5s��N#�8�A4��D����8�iv/x��W�묈�#�^��Ԙ~�)�<`�,�B�����m"4����}��� � �A��$��G>������uN�k9$�HG��Z$l��=��4��)��Yĕ�ao����][�>3Z�~�h����&�N�r��	��x�����#���w�����7�U��^e*���7K%@�Ro4M��S;�z��R��>��]��4��U_�XeSB��,��uM�Bˀ,<�Cu��qBҠA�ԍ����ex�<�v�=�-�2gH��s����TY�4�K�g�C�Q���-�C�_s8=vvX���E�ÿњ�17�3{����Q�S�d"yLt�/#�pRZ�=uӿ LB�UL":��$���D��ajD�N��.G(ѥ�԰&Y�wC�Ty�K�X��jSy�A�oc]��X�Ed��#�>"�*�����c����(�Ç^�J��wB����e[�^��'x,Yޯ
2�O�X$2���!���=	u��G*u��^�uM��^���Z^�jn�;v9s #4�D���lN�N��ϲ'��h�H���ls)���[e����A�:q���m%�I���8����α�S���QŢ�j�	�u���m���Jh�h�S&�H���Yb���Tf3<�ؽ�� ��{e��.�Cg���Gr�Ҁذg0K)�u�������X�vT8���s�U�?��ڐ[V@kr���W���Hm��":�8�7Ԅ�(Pd�u������2m
6KN"��Щ'�S��6R����N��C\�V�@�C�y7���rS�Ř�����k��ʛ)0��R� <R�����9o��X���8�t�&��2���}�Ą��x�UH��m֘)���A)�%x�s�'��pZnU���'�^�g�2Q�ss���(�U�NSz��T '3NU*�4�纱�*���E�������i.YP<<#Bk��1��*|qa��$�8~F:r-�K<���7�E��C�zF�5�������t�������\G�5� ������1ʡ�;�j�P������9B2��?R��n��t��7�N���<*��`�D�+Pw�m&� ����V}�sȩ\o�#f�EU�ЭY�*�K% ���h���X�'#-d���� ��"f�.4Exӕ\�t������A����O�Y��*YMY
NGBCxO�^��#R%.�U/Z����[�yGf�������!�U�m׸AEVY6�H6P�7,)��_�@sO״-�):V�K!Ŋ�<U�i��V0{��< ����ҙ�q`'9��;�
�PZ���đ�V�ѲmטA���C�����;��4{Y��c|o u5PXH�k4䲕�������{AL*���q��˜�G<m�n�0�a����Є�By�����Z�;�xACn!61�Ǹl~�s�L,�`�˰��LjYkI<