��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W��5��C)t<w^��@b�)�aNRw�};��XYI52}��vS�vU�VȜ��h�,3)�$4�7a�-���or(�D��Nć�Mw���tE�N�{*� ��Vȯ�e����D����珗�}�"�m�@���4fS��6�h�D��j�H�x0�2l������b�UБ�ǲ���]�>\�28(�J�V��PᏍW\|&���=^����l��8i$$��z(v~?1Æ� ��md�v�/z��,�>�P� �1%i��Z��H�[��U��G� �����4&��GJ-�x*���d�y�Hg\m��P�wv;n\�Y�,�~��׸7	<�Bt0�I�M,�h�-^IDz�$6�Nԫ�(�\]GU�ƃU.�1�c`˺em�(x�j"��.Eӥ'z�>RӌJ��Ig���U���N�U�n����e�N���Q���8.�?w8Y�)��}�k�����g^4���8����Y������b�5J��_����F�mcXO�n�Rr�����?�W������$d�Ϊޮ[@z�EDU/�<97���e.�^vQx)M݃�t�f��8�T%٢\�_���gu�g�p�Yi­
8��:?k�*ѫ�mn���������T����E�����~�lj��Jp����J\;l�0�g��������,~+�C4�֘��`Ea,C�ͥ��}pǭ[��"���T�pyw�����ڳ���׼�d~3���ze���I}�c��F�`̾P�$V��n ͯ���)k�+?����Ũs�����Mз�)�1������/v�s�d'8����@WC?'�;yMh�f�|�$��k������ݓ�ڜ�"Kt��T�Hc�� �!��͋NNR�%��d
��B���3M�gK�'�P�� �� ��L���>��L>T�UDL�=����<��9��V��ǊҤYA���!eh[~���/��g�Pb ����9�����o�
�����+qu�y�΋'
���?h�Xq�3h$ގ��WP&���M�L9�eD�:�`�V�f��5��Zb.U
y�쓒Q9nkۈ� ���)����:�%!)� �n��dH0���*q��]j����bi�13���T�o���z��F��NB����k���@��a�"i��)Ukڟn����B��(��(g(�T�.�'J9�����W�KN�o[�:���v��|j��]��x
�P-'�*�	n���T�t(�y�Z�$��BNnL���r��
]�����A
����X��\izSi���\|��<G��R�8%���v��U*T��^����"v;��<#[�7ed��E�׸w�Ǡ�Щ�6���E�H#t)��(��#z��5	��f+M��.�x���hz�	�Ö~������n�Nk�'�:�P#+���'d��R�� �x�;QLY�z۸&R��G w 5�K�jh�I���+F�`Z������@�J���-O�����#��8���"��y�{�[=b���!'��iY��2�#{�{PXB�R��
j�nt��'o�<��د�2�|�����#�;���*mW.}!]�h�R)���rd�'K-�X�:\�����v���Xs�1z!�:b�Vu�ZTD�ʫe(�_��Ó����q�6��T�N��Z�;@�L}y�M&��'�l�-���H�M9{:,L�}�u3��샹�jD!�7�oS]`D��_���Y��T�L�	��hx�g�	���Z�����oMt�;H_��.^Sb�_�߯��_�
3'�凝���{��؇��Zˈ�8K��z	u2Tu���9X��Ў�:F�"���ǥ� �ٶG�p��+���>=]��a�`;W�MSz߄�����x\3
(�/y��FȔ�H/Qi��p���ٓ&N�>�#���T��%�@Me�6��#D������x笺k��J���1ft 9��p,���XY�!�����D�ٷ������B�=&��l��h�p�$�m�ڷ��]��YN�ƹH�͙ 	X���w����r�ni���W��ż��~?�w���w�J>9y;p|�U٨�s'ϳNm&����Ȝ�����|ˡ��F�%}&�4�:�uR��+����w������r�{���y�4JV��[�?�>-�j�e���"5[Q�5�V@;�XN��+w��R�Qټ	����M樲zރ�*��I��D	��OF(��Bk��h����O���[n�}g�6��<�țѪ�.���^���U���n��!"���y���Y{��r��Dz�v����	�]4*���>��%�E����_�`�W�����l��D�ޏ�#�x�-L�����#4�����V�[K̸*>�㮙���q?
iqo��>4ＶL�;�k.䭻���Uz�����NQ�Q��'��3�
 ���w�^������؁R�ȇ&���֮��2LJ.N�~�&]'�����+��E7J�0���HV�Ot-�3[T�_$��}q�^��Va�i�0�t��U.�>�2�
"a=x�k���Je��C���W�s+^tU;?U&������	u�F����c�k����9RH�2,e;��A�gZƻ�iXG�a�@|S�uf�[���U�18�ҫk����G�C�$�?F�/6;H�e�7���z�U����b�6��x���e���X������
z9�F���E�@b�����ŧj�H�wS�#�W4L��͢�8���5<�]Ux��gR� ��,8�l��H��3���M�><]&���Tn&�xyz汒`bU<���d��q�߶��_�:��W�5���9����Y}T�`C+�0�D��)��[�%�����C��"@o�����8�T����ن.��#{C���׵l����U�dJ&�����b`��ъ�C8~P�ZD�Ĭx��al�~��0�<�$��	�+�P,��4��8�`��$K�0���CVi~�Ax_�^��+��:J�b
��찫SM�%���o�飷�黇�Z==Z�C<f-Bq�1��Wk���s�ýgu���u���#� Ij�T�Om�n�� �\*v�]"�z�we̙�����V�u���K�����e(��.�;�8Sg�Ź��!I\
���?�[Er���~6;����<@��K�,g����Uy��ݺtMo�2�0�}��̱��[q��S:��9�;dh'��I��EV�Wɥ��Z��9�-:��3#�,1�S�Od�VY���%{����Z���d�<�	e���tn��7�A�h����,ԵBѪt�3H�0���7���4�E�-v\�Z��Z �h�t��}�>����7�W\�	%A2�ngF��&4�3��e�,CJ/R��q
t!��>y������x*���1�\[��h���տh�?�RM+C�-�
X}�և�~%�w̾+f>�bu"l$��'���a:_>Nv�w(�bmϛ������db������%Y��RL��(&~�,���2�q���`XC_ly�]��QX��.&ڻ}oR�Y�
��~W��ir���J�Ҭ�p!�7��T�$2U7
��p�s.�E8��*��W/�)(�{��<����w�H�r�9yu��Ƣ�>��17b�6��[�b���`-<n��m7����������@�w��`F��*c��C�:����#R�a��%���B/�Oim���UdK��pq\���V#�q���[�)����bH{ɋ�\1q@�2\T>�����0O����(��(T9���%�=9uC�Ugs�
l�B�
�����X2{E4sTPQ|��K���C�ۏQw�ϣ�"�*��E�0�K�F��+����������Ic2�����N�UW"j��_�$���i�� �^��IL�����W�ƌ�x��A���z�wx��v09=]v��8�����}�-��H N�Fʾ�+���;��i8�'�<�k鲖3Ֆ3#L��B���1�8���V�������d�4�\��W��pٹ�����8�
H�"�	h���w�?r2��-zUȾ�C�oI�އ�_�t����1����S�Zm� y�E��S��j�BP�jX�H��L�������r���U̒	z�Mgö��T> >�?�VOw�*��"��h���'����&�6�KS����#ɿ.3�򏱼{D�g���t�s����`LeH�e�v��f��M� l�Ӱ�[�fj��q�ʑ����=�� ��M$��pX7������h�!-6��D5.�R��i9 PI��Э�/5��\ͺ����bŃjR��M��h �!�/?���4B<�t�#����;,pT��+|�#�A�J���m �,ʻ��jh���z�T�y��s�sr瘩O��	�0���3�*�lZ�}g�5��甙0��؞)��Ɯ8ǤAіי��~슬n�Z<S#�����.�E{�?Z����4Km㮘��aY<���N��fv�ț1&�dhx�Q��-��N�Ѳ�V1��'v�w�n�A�+1Ƨ7P�i���]�X�w*�s��'�S���ۇ���Xu����~`�0�X�-��ș\4�5�D�e��+���w	r�Z�Z������3��R�
��+ee�nS�) _8�;��p�GW���0=B��oM&"5��{��X�b�}u��D��}_f,��{��Lc�W`����r\���ɶSn<��KAW2R�O"d���պY�WU�K'����yW�����`��3����ԅS��.m�Q�?LFY}ֿ�'կ�7h]��@��нl�l�mH�|4>�x������,\J&�Bg���!pڅ��@f@�Ҿ{Y��Rmu��EE�.t+<U��ѽCo;���Ac�,pA�/֩���l��󀌫|�Xd�`��Ǜ�!V��7��>�C ђ�u�v�q��q/2(�.�<�<I�j�Ի7	�%V��T�u�Dq�D#�{ �ʤ�H��/�
8��fx�W۔���R�E�%�ו֟���eS�=	�4�GΨT�7�k'X�F?�@�2�"W��g��jFL4?�6L�ۃ�|�+�pec�&{7��n�G?qfb�eS�	�Jt�S�>�K>o-�!��i��yR��@�<��R�g�/�Z�;o	�ҷ	;����,Og}>��q�A���3�fr�a�ƛ% M��w:�92D<lٚ[�\��Ք[�\l2d������g���F� �S}��CqlbJN�ֶc��t�K��P0DDλ*;��X1�]�am��,@��(��C��P�?t��B�eN�*�෭/��u>v$��yv��_�T����US�MƓ��|2�[��d��cټ�cc����r!��'��$��˃5��b8m���{�����ڝ½�Y���,c�'c����$�ĕ^��U�����T �Nyy��k޽�P��t��>ݚ{Q�t��Q��h@�����PW8�e�Z�RV���@i��\�e��}�J���s#&�:8�N�AA���l�)܇M�V��W}�yϧ'T9�_zw��Mvp�޶'�x=�����ښ1�ɯ�wTaW����}��9����2?��N�kwl��sI������n�:���b��<��J�d\�Jb�،�rW��!2�N�v#ð�:���s�l���v�-d������[hƇHe����j��\�ik&ނ֪���5�'�=��B.֞:�#�}�E1��u�/!�BC���9k���h��t��N}�ګ�$�R��BO=ǥ��!�S��>!�>V�y������#����v)7X~���Β���x֐+[V�'&׌�3�s�R�a�L~�ܓ�,b��;��O��v�y��abf��'���̪���\R��I�{�!u#[l\#�˵�kZ�x��FJ��,t��z����r�Y��O�3�o�wŰ8Uv�����JG*�ȎT�xg%�����ο���jx�F����I�ڣ1k]4�#�YJ5W�@@̂#=�.�	���1 �J�#I��Oc9ЅNuQ�pC�w����4��+-�z������*���j2�����vӡ>�	��M��5 Zݓ��M����=lã��1�Oa�P��[n,�(����v�W[��,]㨙��Q�_J{½�v�[���n9�{��Z�`}�-w�qn��ҚC ?.߮�]�<iK��޻����%�tn�����]5Xw�E�����V8�5�t�߾�O��|3ށ$���%�C?������]�����
,0��q�P*���-35�y���.s�M1\�����I���x��Jf)��b�/���9_vj]���p��F�`�.�j�e���u�JC����е2�0�McZ���c4�R �6:VFa/�� ��d7�Qu�bwἷ0�,���M*�X�~c/U�P��P�VJ9�(�Ve��g�5vLV�I����YM�pf4HG{��k�,����Bƶ&E�m���x�S'�%-,G�P��Bvg�sUeM�\�eɍt��#���V�cTj`83�s���mlօ��h9@b�{�ޥ���e!!���N�����Y��2�u�}���O����JO��*n\����T/�����h����4Z"_�I�iK���L1j��I<��i����P�u�
hA4�u.g��-PL��4�eG�x�R˔����"�S������k�w j��0�K����ו��Qе_�V�t��8US�� �=�v"�+������_�k�no�x�lb����q�f�5Y��p����G�����{�皿�V�s'�W7��=��S?	
�ݍ�጑��5b�W
f�A�� �h��T�]A�=>�c�����/aK������l����씞���ߨ��h��-?>�*E�^�~3�-�98[r�!�������[�̘�䧌�D��V����D�Ö��U�����TCPk��c)l�6�-JOF�&$_Q����u2�ؖ枵	��ۂ�񏔳�4\�j�6i���d��S89�Y��*�:��" 8(��4?:�nm�#'��~�ڄ�|߼�Z��瘍��n̍CǄeб���;�h6�Z{��lS�+��E\_��- K�14ҷ�S�L���[Q��D��w̓�h��\�cؐcQ:`�b��Ån�ҳ�7�Ce�S��!a��/$��^+�m}�ǈ��8I��~�Zd�����QP�ӆ����B!�#Ykx�k��TG�o�8t�i<�`�Ăm���Ym����L`��+~x���Z���F���q��-*��3p8�8"<�ሜ��,ۜ�)(91f���7ņ���9+�Qva��A�TF�v��G3��xBl�ʂ���̼�z��,�(���]u5�7|z��ɋ+0氍
���޺ ��!k�f�Q�fգ���|I`�O�x6�,b~��Ϳw�kmĶ$��a$	,����;a�9���X�f'��F=�#��i����*`]�?����Ӡ�j�0�.���|.%����d3.b>�`b5�<��4狘/�ǟS~�%���b0��L@�h`��&���T
�
�\(NDQ�u�.+H�p;�<��
<xݨ�/?w;��������JD{��Խ�|����"tY��?����;��n��_8CH����C�]�����I�%���H��`�
E��"k�$9h��]�,zh��!A�l��ٿ�%���^ٗ'\��h�:����6>W~�<�X�x0�7�:�y�ͩ�C�37_w+�d�r�6�"����S�Ռ��<1�i���1
)ȕ����S���I��2��K�|�VuPf�H��}FykO��{h��%�g����XZ�ux��CLh��B���^���Y^u{E\�y�gP��=����g�P��}��V�jPw26&��S�S����:�E�2]|�8o���y���?�����`�������6�Jh䳇��c�CV��H�>&�$n/٠��W���X#5�.����Υ��[O�K�h�x�{���hB�!Hjfta�Ze����U�c�@��M�w� Jy�$~�<#Q��H���<.o?��NP��')Q�~����dr�J�P���ځ�s�'�e�G`6{p˸*V������z3o��xجQ$u")���Y�}p3�ۇ�����#7��.�׀���-�K�ھfU�2ߞ��c{zw�/����̑�p1��x*��������R<��)�L���86�:�i� do�u9J�ߩ�Gџ����S�zT�4�5v6���H���v-A>=�����HXK{Zw�tu�Bz*����"�@�&�86�����(Oi�t u�-�Lk�YlN�Z̯��I�E��C_�Y�R���)�X��O�O٩��0>3�B��F��'��E᫿_c��A-���r��ǲ�� ����~�G��ĩق���Y'��X�h�P��uj@�1�ln���np�&��޸D���&����~�M|�Br��b8 vq�+�@���n1��|6X^�r�MIz�v�멙k]pJ���%T�-�	i��¶�*2�{���0��a��/�~77��3\xM:�-�s�|t�
��(�[����(�<�c���s���
be�e[�@`����>��o8�6�ҹG��J��.�1ky3�Y�n��)����Y��蘣Q��4�\P�~�_�%n_� ��ePa�E0:� �:��N�������,�����F����r�Z7�o�#���j��*eP�c�	�B�� �x Ϯ���d��y�p>b��8e��󩐈��a����ނ �y�A�iE��1ؼ�(��m��O�L����X\3���B઺�O	>�ʙ#��!  #�N?8��/i$=x^(�2r��3�qA����K��|ɔ�O9��bNG�M}�:+��'�:�""�4Q6NUp��C�dk.!�z���G\Ǣ�S�(4P\ĉ��q����W�����hrj�PM�^��������>y;)}n�BN!�/8 �~�	�E�ȟN�V��J�SҘ��f�:x�4��J�������yY�����B�B>i��^L���L&�����3s�]E������=���7�m�3��N�^��y^�����(cf�y���A��{o �N�eMb62Ku�o�-sG�����~_��w�f^���74��T[�2<��yPG�}+�b�D�//���h��A�_?�CvFdu%x��F; B�J(Ґ�.�GZDZۙ�.N%��{�d�ɀ�{�J�iJ���Q�h�	����_P��\���ޛsK6��Nu��Sή�A�q��J�( �¬ǈ��H�����M)Z���^ʢ@w��A<#.�{�lX@e̀1^��F�s�h9B�uJ/Ɨ��!�z��ַ�u�<��Ђ>����z!��Q�D�\�~	Z��4 +��ˁ`�NwŻ�kM��Ilf}��0Y��es=E�c��;������� �6��
:;l@L���'I��Mf3��X���e��	n����eu��#;�pV���t��"���zF��۷��b��om��.�7r�Լ)܀_
�f�*�c8��<�$�Ң'�Q���jM@���+�����,~[U�?+�$qYp�	��'���z�~֮S鈗����� ��T훪��m�_f�t�n:f��]�]}6+tQ���������g=�SaHM���r\��V�=tJI9h������x��{u��W7��]��T�/���~�vk9|���<sī⿧�$��w��`�ш֒U��/~r2�ro"G�h�-����3Æ��ԝ�[8#c�m���k�Wb����zO7���´Iw~���ThP��Wr!'�dޱ����N�X�ځ��Or�S��\��(;j��h�b?`�ೈ��?��EW�Xe��v�L��b�6៭��/]����OK������,�����<�����U^���v�����_-���+������뭩m��Y�5u��)�UT�0�G����Q)J�.�Dt�}�~��4�w��ΠMl���`�JDB�͝���t"��q����Pk���`�%�6G�|���b�4&
*=~��h:L0���؏���g��\�*�Ow4XIC��r�h�?l �iF�
t�2	�?#yI�W&rax��kj��s]���6B��
C��<���{z�2��'���S%
��~�����|���\\����Yad&{&�d�ć���c��Y��U�Dև�Gv�T�!���(�u:���q�.џ]S!���8�ysp���n����6�Q��(L��kp��ov;�4�����K�9����v���S;�aIB�x!*�TP����� �ܫ�gr�?4�,(�_�\2Ag�]K�%Re�p�����>�t)����U�mH���է�}3�P7��"�@�C~��-�����w�A�#a҉ۂ�������*}/��ez�s2�M<�(S�u�����F���`���yϗ�q��ND�w&*�#4�4��G2���l\ȵ�2f$\xxFS��kފ��F���Z�D�1i���g �V�e�����\7�6����զW���)�Z&�) H�.}���W�ѿ�_����`����τ�}p�P�$�b?_	�����9���4��A4-S�����{j�O������ݤ8iN�6���iޘV��-�&���9�� ��_�N�1w�U�3�����u�To�<JoQ��Z ��Z9����^��x����[�3�̏.�������6�~�Ӕ���Gt)�W`��ø��'7*m��ΰ�؂��@Ac�Q@:�4���&�K�1�F��/*�<${9�����ZqPJT7�k���N��|��"�E����Ou��@�a}X��Q;� �L�QwP_I�Q�r�Ѕ�ԍ��.i�Ռ�눝��o��}���Ѡ7D\�W�C��_��S}A7m���72��Y���SJ)�ݑ�5e�K�aN��T��XzDtكr��+Ή��7+>�(�v���������$3�K ��f`��s�J��-�"XY"�':�ш��	��.(6�X��P�U�r�v��Y�;����5��f_'��b�-J�џ�򖩊�C8��(�E�hԅp�
�8��{�D�0�8��Êb�R<�����ovSXU��p��'���kn���ASg�*�1m��e`W���IǗq>�kNq�5ssFL�	9�@A���$=5��>����ߍg�#�3`Tc^����;��ҬwGԶ��~��Ӹp��f��3	F%��Jَ�q����|*f&�	st ����E�J׽
�Ξs�}eb��Pż���k�7 ��=�PS�tLd��&w1F�62RGܗ�B�4�����U�������	�Inl
 R��@^��fƂ0������YiB����4��w�b��ܤ�����轡�������F�-ϰ(2����R�e$�f�R� ��ڭs�Wלn~j�vKsjN=���릨�:)C�	���J��IQ�hbB�"�[�~�����'��(~}q0H
ߠ�	�^ e��`B��$!m���>�>r{4X���[�m_�7�oV��,gO6t���d�m/��b4k�e��+�2�*�qo*!�܂�d�qRK�z����0q���u�EI0���m���|�e�y*��FJ�WZb��¤�@#��%��!�����e���m�q}�q�Z^��N�C:������Q�:���M���F֑�4*B�Vp(�}���9i�����}L�/�l1!���sE]��e�#cݧb]��[���u�����y���%_�g��V3zf�Ь(��I�(s��X��ȋ���ƅY����U*\�[ۨ"K)r�c�Q~�k��5����V��ܧ3���ˋ�CCZȇ1�i���]e�W�ص9�3T¬�*�0e��;�e�w�LE�R��%x+~I�KtXp���Y�4���i���rnї���v�y�X��#�[��JtIM�F������]��"�騍U}� �H$eT~ط'_K)`?��٩��`��j�Q�+�#�X�'��;�G��KS��x�g��}��ɸ?VA"��w��+6���V#������3(�P�疐6�ן9r�?Hd�;X��P��1K�������1ν�%�J�"@��!�W�{D̗�O�+便O*��;[G���v�|&|yD��p�����g�&�J>��ԣ2oS������KC���%#�%|q~�|�s�ç��UA��-��S�0ig� �l֮������7v��h��kK�O
Z6�c�3�~^� ����n�_���!�L�Dwܫ�T�猜������1S����~�)䚽]8��P��67�ύ�u��E��V]S�	?��nr����z�1���'"'1Cc�6�_����������mqs`b�]X:ϼ	�d�k��GXq���N��RP5��8w�VO��QK��0"��X���"��c6���M�9�r�l�Ɓ��
���4��Uu�1�=x<�0�ܟB�ʑ���@����x��d�$+Jj/R�R��1������37F=�������f(��M���@��SNs[��}�t#�
�yJN$��B=���Y��Q�q�&m'�o�[���G!����a^�nc���붢�� {�n� �P�b#k1y�p��@��ɀ�a�u	�p�^�����FN���!�[��)�߷�@��J�3�ۖ��):��7�{��w{*�n�@K�xm<H�XYR�=h�Bb�vz~L����Y`Q}W�gˍ`lA��r�*�%��]��Z��AO�+�͋B�U��&�+e���s���Zg9z�������Cm������}d�rO�M����+=ƻ%�9�{z�"�A��Eݨ66Vzt����-51����E�I��r�1�K�@����=�0��M���!rQ� �ۡ�wK"���`׌G�F�˃zF*�3�y�*�(9Tb��@�j���!�W��8���k�E�>UX���FQ�m�X���?���~��!�y��`�=�xU����R���H����+e�>�H�G��T��˧*a�Q/r��a(���F��ɞ���=���E?>�u%JC��X4]m�XI�~3�(�����=+d���	�ŐJ�D��t4��[�t��K�ɳj>��hn��c�O�"&/C����ك.��;,X�k�p�a�1� g��B�_
�ܿeA���R�r���w�:�i)�'�(o��:�^��<}x�>X�3Z.�M� �'�	y�C�8S�3��t���8D`��t�SQ&?j1PCb�'({9U���9'X���BU�:��UDeq�<�wT��B
�2%N�����ӷ�x�FBƅ�G�� }�i���8�j�(�n�*OX�=�an�#�Cˋ�ʘvN+�W���yN����V敕+9�3}Õ޺����vd�������R�Mr���!�8/�b{PC����]�#�_~�=�z��N�#m�T��U��T�Ȫ�q�.��s�y��o����ӸEK��wC|\J�汈OSP�П�nL$W��y	n���\u�����Ȃm+���B��ws�n1�߈_�v���\��S�Ku�X���ǅ��
%�)�����=tH� X��.Tb��A�����`�0��A����̊N|�t������O�pɥ�,�3���>H����R]���wD�;����1���|<�W��*$��}:l~�*es����DT�!��t��`�
����ۖ;�0���4��OPX5t>�6�\rɄ~�O��FO�fVڪD(���*�������AJ��s����S��n8:�_���嵊$�F��p�,��I��b��F2_�G]���>J�\H
'd'
��a���?��m�ގ'��v懼:�,���2 ^��i޵pPj,�t�w�5�/nt \��^�6��KVk�;����]���D!�����,��Ό�.?Y^g�t�����e%�r���GD�VU�u.�s�;�F8|w�ʰ��J?�񔘱��+�`NM���Z�dM�{��8|���6�G�`,H��-�V�)4y�0��Y�f[��8�x+1���D7�L�^���1���w�J�{֦{0W�N�M��6���bK�0���0�p5��ɿ����g+IQI~x0���:�J�n���s0ἡ�İ(����P�8���;�}{'���4�B���}�ri����Z5�i��8X�0�QWc��u��S�ɏ8�)��iJ7>=Uy7e�	���6o?( t�� �~���fu�ÙV�S��m>B2:��j[��+�X��z`;��ȋ�hN�����j�_}�n�>Ě�Ӯ
JB�$Z�c����j|E�#��قˀ?f�e��W�|A�B����>^�$���<Q�q톇Va�7�񥇸(C��wǖ������1m�}+��1���c�"��=��j��8݅�j}`<�:m���ёO`"\Q00v��>N������X烧����1\�}K��e������gI�lb6��Y��#K����ا�<c����Ҍþ�_�P�ჺ���l�Z|��9��枯��s�0�^�t�X�:ߏN��49v�$]��)��v0���Rȋ�X���A<�Ka_�����n׺��������;Z�'9͌�;� F')]l�����Y�M/�˥�A��)��FV��fv�}b�YS� R��ۅ?b��r\�9�l��ɝ����9��<l�8H-iNe���B�'�+�>�t��;=r��t��q��8^��SfR�՘]m��@�|�ϙ���G��̛�Sh���y�Lzˆ��$Ǧ���+�#'F<X��G�@�7��'C�	��Ǻ�;���sWpT��br�9���hH�s�"Hq���p��k��A�7�AC3O$��َ�h_�������*R�,�wrI�(��j�)��5���p��?��� �,:p�r�K1��}��MP>9nw�O_dr�pn��3��#g:>r�;�-PfrG.��͢&�4e��U�1ט\���d����'!z�B�h�o�|
�េ;V��)��˃����AkB!�����59	���R�ھ�osh�.A��u�V�4M6�������O�_�ԥNh`��ʡ��/bA�	 �w��b�R>64�ܚ�u���}c��)͔�s�]�!
��i��c����a����G7fGÌ������f���
�O~ ܡ��%"eɖ8}����h�ر�e�������8�UAC�?P���q��2@>�UY�!l.eʉ_�w�}:�P8��זO����#u��Hv�N���8�?�~�hU��[;Z)~��.S��>q���8]b���)��t!?�����K}�mѺ5��Z_��;�2Iͺy�P��NL~������DϋNd��bLC�F�k@\T�;�}5/���z��f��j�P-5���@�%��1Y�I�N<�	��_�f�!�w�0�Z�I&���讶v�>CH��� Y�ĸ�T�.�}�F�G9����������`~�)d��m�k�/z��"��9p��wc�K��90�#"ģKc�h!���·m�z]h����8�c?��ݚ��w}��Na���"ު^����oE�e &�ߡJ�����G�
���v��up�)�Q�R�dMK:�`L�8l��?R�l��b����Z��Es�dnKe�n��}oz�jr#�
��q��Y�`��ciCi���8�,\X�*b�1�������vO�Z�Vّ�e��!����_1���ED�[e{v5�&�E��>ru8Z�ؽؖ��h}���8G�;\x�x6�h}�Į~���#QHAf�Z], ��w��;,xiƼ0K�m+A���o�����F�S&����8��cY����*[K����5�֚�l����、�>`����x���o��R��U�]1ӫ����JƎY�i���>;9�x(͡AZ�ܻ*YG�%E���;��޽�q�^�ܳ���+`�tmc��u;�)��`�=��>[����)D��X)?��3��O��@��&+�����i�M8/U�H�#*���6�(%��Dc�xƬ'y�K�2�_܋�i+i�5N�ɉ����~㜪{K����Tppg��g�A�j��D�	r��w �r�~�-t�C e�8
�/a������=�}��v�I@l20�k��1>�R�i�ʕr���\D��h�<E����	�|�
po��/��D���=�޸T裼�d�Vk�K��Iο������F|��B�#g�q�D�o{�Vw����y1���W����"�΅��U�HH���q:����j�ʧ؅oa +Ն�&��E`Avz��v0��J�}�=��5�Du���?���#�sE%��a�\O=a$oy�b��q�r���%�	�������28:�i>Zf�; W��VО	�MLA����bC �.�B�:�<}@�W$_b�����:�#ťh����&����P[(�_%w������*��iB ����k}Q61zyY� ���y�-k7q?Ԏ�\Y�y��H�dc�(��ؑa��c������Ǖ-�qEL�{��T)���:ɟ|��	��R�HCZ�&{�_�iѧ�[����˜�\�zvQPЕ�c3n��~�Iwl�����`�@�`���>��T�{,��� %�?�	�Қ����?�mD���^n`W�y�����JE\mP�ξ�`���?F�dpa����%w�in��~�6�:ў~ϟ��g�Y_'��>�Gag�O8|�H��c���(C	s��pb̲���U2��6%i�혳Dc�P��!���X��G���B���n��w��SXh&.���>��*iv�G^�~S����R&#ɜ5y#�����ا��XIH�w�1'�M�'n����Y������'�K�m��%��c�l����\m�tp�dXK�qׇ��L5�l.7��|Jة��S���H�˄p�;��m��$z����ƅ��C�}��Q��޷��Nt.t�X����\wo�O��n�nmI��l��Uz\���"j`���/Lv�ÐUtn<o��X�+�|�=~�NO��
�3Or)L:�p�$·\���L��e��$�Wf�s;;�K�1���хNi9�֞6X�6�M]��=1�I�[�a�LƤ5!@����f�1)��I	�L���f�
�.�1v�р�O%��<gf����B��J-���P!�����\;�ϫ<���"��L�����r$�2�*e��Zه�uJs[Y���J��{���h�x��ii"�xO���G��bgf�T�����i�cl-j�(���pڰ�6��W���j�H%��R��4)9T��_�A/o�f�{�溄�� Θ��T@�t�������>��Ԗ���t�P���BؚUo*�	 (>k[�`�V�A���A�vkM���p�P�j���h��fX��Dd� ��~b��5Җ�wT�.�����\:��x�sV��	*�+����m����P9�Q��26I�R�+DX	�Iz�m.�<�П:j[����x�h�D��ى��n ��~b�����^�GbS%�l��J��x��h�Z.Y�(����+NdG�.!�:���
�����o���#V�*����c?㨼����`[�fP7�#��r.��_��.��r�����<E��H'~��R[�a���E������n�عą�c�牷�7��{z��˅�2,+�a�����"|b�Q����O��e��
��_P�桲Ay��ո�d�3@�A�L3�T��V��>6Ը��lZ���@a���mbm�%�a�:'���Y���̢aF��-Q�5�G��.�P8��W~d���lQ"Uy�{-����C���'�0%˟Ǫ�+��~���9��rB�����2�����)v^�tw�܀�"�WSl��i�QB��������*�}�;E�(�X/��^'��8ijE�\���8T��y��n8�,�(�����4?֛Y�X�@���6a��c;ۺ$�[�+���2�/���8q�
 $��0�5�x�o�;�J�%�}"�'�w.(oT�*
�&�H����`�:#:}�3Z�����,߶@�5R�~�YLN�2��NҼm�zdǒ��؃]��Ѽ� %b�z;z$��,���ϹH�V���*<�dVNΊ����f�)��"�R\A�ɫ�]���d����c��m	��Gn�;��%f$���8R��}�ޗG���f��%����C��+��\������y�~��%��JYGb�դk��Wd,��lԃ`L�UF�+�*� �{b��d�!:�Y�F=3s�hB�z���������b�����!e՝��ci�V(T�s����9��}�O�>��2f�G$J@%��j������^���p��+�"����(��8A�Г��*Zu� ��;_��&$�/��/�y�����'����!�B�1����A_���p}ŵ�Κ��|S�KTt:��3�˸fJM���3ER���y>�IZ9�6�5����^���yA�����~�n54�\�
1
1��h��d�E��Q������ۇ���t�ۂ��+O�V<o���V��bv�'��4s��6{�D���V��>������)q|��l
�]�S�St35�ƁeM�Lt���޵n&��u�O�E�=)�31�fgv��;?�ҥJ��̥]eR6�~)��,�=emCÉ�Y����K�f�*��r�h��)�������Q�/1�p�z'Ӥ���HI�u�˞�JƧ!��s�����,Ճ��t��O4@\�������kM�17��1#�6�iF'�Ő };�3�}����j�uZ��'zMh^������HգZ�[T����]&����~���xss���!Fe��@+�gyy\,I�.1�a���?���5�(�u5�ԧU�w�o�r@ڌ�<'�j��[���M6� �����AϺ� h��s&J[d�Z�>���HJ#@��#\p*�3�#L���*Ƹc���MKF�:�_ơ|!�n�Vk�X�1�DF��<Z�g�^�.@V�
H��P	v2��'%�0�����E_��GB���CJ�x�\�a�'�bq#����%Y�o���]��^���U�W�߳d��c�_s�͌m��T��2M$�h�Q1��Qi�h:�<_�ѧ5��fk��IL�"]Zp����ȵ�Y9(�y�C-�@���D���8����'P�[`���؉����?�� �to�5m:$3�����7�!��q�������Rk��n�atǹ�V�^����]���nu���Y����͠j(t+�Qs�pF�������&&�l,r�$�
y�*��p�j�5;�� � 7��^�ɝ������*����?
@�{�ĺZ%��J�~i��}Ξ�
����"��Y$K�e�ca�ax9Ǣ�s���k�w����a������2�p
�Q���"���W�y����i�͟�znE�;��)/�ߙ��1��{��X�c
�Z��]��/oJ�[�80.0��	����d�H�@(��R⸓�^��L��_�/E��*)�Rw��'|͑�^2��ӂ����τ~a5Ճ���Y'�v��P/R/ϔ�0>y�ɸhHV5��w,^�иk�57�L.h$��h�L���$�#2 H�Y���TC1����L�7�a�yi	ݱ`�l޶ӝ�zMN���zpZ_����oUWQ��7/DFlN%�����������32����T*T��wb��[�w���ìQ��M���m7X-�F�n���~�Y2����j�?��T���T/������֒`����\�}{w��?��7`�Ih����)�]�ǂ�~dgBơ�cQ�Y�%g�栠���/_;v��lq����!`�:W(��������/�A�;W���G�q1F=�gj�U=���ûC��,�By�L\- ŗ�A���z��H�3ަl~��Y r-S ��MPF�>O�"+5e���[rm6�Y%��B�酣=�\�?�v��b������ՏsfW`LE��w�O^���A��S^����>�][��}ߓ�/�m�cȮ�	_{�e٫�#5��>��=����E�dC`�{?�.��D�(Z�PkE���"�,����oMc�;@s3./9]&���দ�ɰ�}w���v-󾵁i ���Q�/�5��ɛPҋj,E�w<�$�=kf��.t��D������U�n���D-_�cn�b��f���swW���z��,CН$7�����OͧP'��� ��̲:�Df��C�x��t�,'k~�Ц����)�&����5A֥�¼���]斏3&�?�Y��V��q`��Y�Ĵ�!�&H���J��@�~	�<t.շ��_oi	Ar���V���d�J��5�]W�Gi[.ǃ&�_Z8�GiE�'�ѿ�#��ڲ-@�}X�)����&�:�e��פu�%�i{��@hn��|v��X�K��J!<gn`u	����G*� B��U��|�^�8A�:�Ŵ�q^���8���=h�;O'�X��UU�,��ox��@؅쇃�i�#������p4���>�s��?nZI��G���>�)@zW^�/���a#N�x贩�|��M�E���zsL�jA�o��r8��Y򊿳��F�d$�o�son���&@tu��������8&5��f�p��.I�Zn �� o���6#�i�Qx��& mu�gH>[�c�U�(!�G�[�n�-�1Aq������c������cL�W ���a�,�`� �M	��yL����P��b���A������*[��gD)�ˮ_��Q[H�*�V�3p�{�-���S��3�*gQ��:��0A�i��pS�ӓ�L�j�& ]�Ď�lk1�%��攅bs��f����?�פ�`:OE:��ܨ;t'ZH��)�h��t��?�Z��?��8j2�J�֠�9q���UM���L�k��Vرˈ k��Y'�
P��+��N�+$���&Ty�����i�G�PQ�E)���@~/�yZ��`'�Q/?#%P�[��:��Uy�W�[J���X/P���1��#|��֊xB�ȗ�
��}�C��j�l��|.)�G�Uȵ*��E��^���]���ܬ"�\IK�	����Y��wF§LQ�6���LȤ��<�J\{��@��lt�=i��6ǅ�B,ک�7�,�"�-i�}����lb��$�!�֎K��P�2��"���h+�5n &Ô�2���"���~�/ӿ�1�C�as`��Zg���ow�3����AI�;}�z��{�1�t����--�uhR�E�gJ]'��7G��(� �ȓ%3���&/IF�?`dX������֕��D�0��e����Np�pS%y΋O@����7Sl1�O"U�VXl���#�0h�腧�d�N�����~��,� ���+ޖ�Kxc<o$��Rq�8�b���]��
G��-o�����{A�o�e;�ֆX��u���`6��/��If`c&nP;2����M�Ȅ�\�]�o�s*�#n���u|��#�k��O�<��e�>�����5h�(>%4]I���N��,n����$+�4a��;������`��|-�b3x`-�.�Q[����p{�=�>J��Ձc���B@���W��� ����+Blr'V��ڦ�1n�T-v��҈��&"�� 2�PReitx|GBL���0�N�0!a�H�/�Q���>��->��ݯ7`I�uңV���`"R����fX��^�j'{���A�?�3�5�~�J�팜]�e`h��O��(`C<�0xUzʣ^�y>�Zd�3������=��p��KKMG��g?gg���H�U��,Tޫ���k�U%Hx� 1� ���t�-Jy�o �X�;�˃Ëg��D��$}��:\i����{؇JV�h7I��Iqr3�
O8Nl�q�-o�R�o�Fd���9
�F�}FIT|B�@��2O�@Q����)*�:A��EbOS&��MSw>C����ېv�蓮qD�W�����0��i�Ƈxu{�X�
�WQw���ds��w����m蚤�ᕁC3��K��ƞ��1�\��3G�����
 ���+3pG���8e��^�%��_K��ɐ{�gp�p$�~��>�%�l3zz
J��W[�~���Tb�8���}��R��k�����y�\I@�B�DڹI�:�����ēHu�\�����刣��o�Di��!�M�?�i����ƤBzbU���&)�Y�F�2?w�2��u��=�;�ڔ� tG����83�x����t�^+_%���2��W�h27ћ��ev5�KQ4)�h�� �^����h��21\��}�D�|�Kں�p ��L�Ԕ��E��L��⥛w���1���	p�Uz�F�M��"YG'	xn���+��K���ShţRU@�n�PQ��q��U�c�!)��^'az�Ao��F�FV��6X��r0�=�}�j\{c�tI���ڹ��@��žfO艫_lk�Թ%@fbF��@r���h'���r��9fDX+�XAa�&FDB'n9�Z�ֲ;�9 a'�x�Y�q�
��M�E�t
�WS~pr��1��y��E�!�J=���n��[�jt�6�U����	���:H�P*)�2Kh�+�9�����k%mj:]S�-d�P�J�Rθ���0���9*��cXGZ��H��c ��H;�`��V��u\X�;�J'�1��CĜ�l����V��LW#F�� 4�A���S����>0�1Ry�u��e��r��Q�a�/`��3oh���:�D)�����V���Bn���us?��\ӂΔ���C0<���$�'�̼�&X+"��3�Q{�@S�kH�:L6'�ȸ)��v�y�v	h�1��@W8��ͅ!�7X)��#��Ń2���=h�&�#�'�����`?�[�N�=9��>������, ����� ��� �Ѭ�	�o:H"I�t����rrx�5���jqX����/�6�lZ?`nIG�Ȼ��B�>Q�д|����5���7��z{�V}J���kvӸ'"����-�y/��E�Mc���/��c2�2�̒���>44t��$�^��Ѧ"K�p���<&!�P辞F�%�����E�h�^��2;
H�Ms�b� �@-
��qC���9ta�Δ���0��(�@/x$NXL�����9G� -���goz��kR�'���br�ur�y1��l�߈��R���M����z��<�UL�|	��#�}9�3���D[^b�{��Eҭ(`�*OG�v�D}IC�^�f��u8�er)��%�>�'��B�0�Gw�m~�%e�
�8�h�Sa�x%����t�5�z;��"�巈��%�0d�"K�ު?��6G��u$�w�6`�?@���"?��z�9�o�6� n�E�� -�֛�� ��j�����.Z����e��O��� Q�w/�.׆|K ��8���b�q�Z���c4w��A	��䅟��K����%�ZB�@�ឧ��w�#_��>>	��4۸P��bf`��,��D\v��Ӏ'
�:��xx���^=C0����렒��������@�A��Sr�M?����;�~�7)�[���#��e>�<f�8�]*�:��#�&�B�T�L���̺�� h���$���̺�=Ԁ���_���>�£�@�����Ab��9v�M$�p02��q�8��$&��V��{[�$���w���s]P�_�rD��h���g��
|���M�W�1��#o}C�&>Z�Y��謬c�����*��]{\cM������17O�����[%�.)�ԁOT��gU.���W��&�V�u�L}P�:���0�E����{�گx]��$�=.�M5�;[Oӵ����n�vS�����}�8�C��.+A��3kJ.'
3�J�/�q��G�N@�C"��Y�ݙ���m�� s2���Ҿ"�����CM|���5 kˉ:�r�^��Y�	�hli~zv~������#|��o. �!�𧧐�l�Z^e����F�e�j�s  ��V6�
@��~U���$��/�NڛmOTL��M�Ph�@�k���	��Lң�i�<��?Bpⵥ3U��$�ob��8�C�zA�o&(��q�}c�@�9�V��LE�J��d�v9�����c�,�����05rz����Y>�9-�A�Ti#-񾟔�V���A�<K/"_������[i}]�ylX
�]6�0�q8GD�Q^�MQuUk�[�h[�1T�Q��δ�YR�B�op�c�����T&[Ү~~o�l$�P��yI(w����w��Ze?H������M1���"����"�[T��jj�����Q�:��<ٱS���f�x���A�k�(���\���+�ΛUj�>�vj���K���L;�c��{	T$���?��SuI� �*@cRe�}��ͧ�b���s���dD��3�D�c5B`�@���cm*	|5���w�: �������hJ����>��$/�)j5���"Ǖ�-Qu����&�_�d�qgf���f�I'~A =�|���Z�S��j�X��n\�*O��6eN���j�V"�,�`��|?�>�x*��	- !��^̆D����u�9��W� ����q�'7�۟��ܿ�D;!�ZH%���%��G�c
G��s7��C21���tX�.��f�ģU&%$8P��f9IbbQ��5�j��� 0�c��+��{�X9?�ބ�z�O`�?���N��H`JLY�)���D���^����D`」�t�	Hz��f�(ۧ��D��������w>�τЫ0�6��z0:�(�M�P�)Z'���zh�Pq�-,�=
�L(�'t������Vl�;I-5��,/�'��^3�{���e0�E�\aBl7�ڢ(�s�Ų6�)�,��7V��	�[��K��<��BH�\k�'�ULrͥƂ�d�*)��p��jp�΍P椃��փCo��s�Q��g��R��3B�$J� �����lVLzO+�����K����_��h�I�"^>Iy?@(��d��<��<>�E�2B�d�c���b�5�-�uh_۠�x��r�c[��q!��}����/W�uթm��H�����@�.���l�"߁�L��Y����	���Ic� ն�I����;D,6������o0���&� �^����9�j���n2ÚI`��b~�_��L�ۦ��ϧ�!n�)���s5ϛ:��ʋ�ᎧLG�g�p=6A���+-b����}���vI'iY��}|}_1��q���B�1�ؙ�s/2w=_�$k�U=u�����c�|�:�%T��Θ�>\rd�[��O�����p�2����o���u�]�&����p5JJ`B�j|�' z=�=�B��i:�L�:�T���ߘ��z�ݘ�:���،a�+����H� Vf��P����Q�˶����r��f�\�M�[�Sw��w����h٦�XPa��`�|��3$�RAL��V�2ȱn��K�[��l��	��X�l�V(��v���ڨ���Ya@�ӣ�t��5Q�j/Y3���g����X��`�ۤ���#*_@U,� M����1�N:߬���Q�<���+r(O����=�v���\w&�}ж|�EMP��X\���eر�#d��oy
"&Bas��>����
�bh�`������ҫL��{*{���^���AL��x(����}]/�uE�ʰ�ؗ%H*���s��E�
�!���Ӄ��:���*b����:�ΐ��q��{ �t)LP��(���.�!�|'a�/�¡�F�q��'�-�B�f���,9|mN�%k�bo=B�F׵�^�����𑴤L�����V��#�O����,͊��2kM��Tb�������78�ae|�H ��$�K-s�Oy��CF'@'	�;m�K�,��e�a܇p���փ>�����q��rs6%�3�K���s�%�w���2?
�'��:�%dB����Y�(�ߨ�� �2߰���W�A�����N�h��ú�RҴ��3�)�K�]8��U	WK�|�]M,�$��oun*//&�ɽ&�WFyE����z0�v�^ES�ڿwlܣBpA�+K���*Z��m8��Cik��a�׊c�`�l�,�.����[���V���"�(�yn�.?uv��Y�N�P��=*Cn�%�o�a�M��-^�cB�qS�^���8��$��r�`��>e/�y�O��ì3�!m؀u�b�m�&�n�6��BZ��:���x�7���3�-:��XbN=�N����	����1���� ��M���<8�L��4\IDi��#E5�YY�⼂b�5�Ou�/�^�X+k�P���}�ߒxl������IٝXhЂ#8)y�be�c�H�M���,�j#�E��k�f��N���Y�O0A��Ȓ�rr�7��**�� ��/IL�m�2�UymFzPF���SmgT�-�#�u���W��8[q�\f@4���J���o�X��Wg����=j�8K�@����"3z�/���P�v��!��XRF�F�l��Yغ�0dԍ�K^�Z,l��p���9Q�)�""+[���N���4K�c�z�p�/7�^J��uy?������mT����Ѓ��ދŲ,�xUw��O���n�7��ix�5tXp��M*�h_��rKR0aj]0�@���{v�̮09}����{���Os�Y3���P��?�k���p-�0��wI�����ѿ��N"��u�p���qծ*Ӕ�A5��+`-���&��%�
��nd�����������US�f�i��H&̖��l�A:�,Z� �;`���B��R��w������)q`ϻ�!���z������1�u"w��-��(��q[������/���#s��m�e�I�g�.��A޷�����6 N�9���S�F�$|'�FU��E�KB����F�t�
�UY��Ӥ�n,��5A��;�ӑ����6hp��R���h�zQ��陓�I���7F�굷��`�{������[|�%m����ȼt|q��$�(�	�s���TB�"�\�k�J�C"�&�
6��)1��"Y��ʏ��;��-��m{��$G��cx�}Bۊ	4�9�]�K^d^���v(E����t�PU���H���1I=@:.��r�w���:����TrgL�5+�lP�� �K�^1���Z�[�ŀX�bX���;Br&�8S<vu��]�mlAO8ZC�ϖ�o����^���t�\���ٸ.����fC��=��@
]m"nA\8��a���k�}|�M̧�8��Ǔ�L �'H��|�G�iz��X��3.���ͻF���S2'9\��%J�"��;\Hz��N���X�Y�$+��P�`D��u��ц�Tæ�nւ����@)�|����AL����t�K��]�tf<� �o�4p��V�#�Ǖ~P�CwleD����Y�J��, �SW�)�N¢���ػ
����&ڹ4a�"��L�~��~l�v�x:�e��i�����S}�-*���mح�[W�ŷ�[�:��ҁF�`���ޭ��&�"O��`0���D<�O�F�`&�#�%�0V��bX����ɕA�[z:=- 0D��&4��#R�q��6�?��һ�G���fŎ9Z'�xBS��h�E�5���r��$�ҹ�u�Z.0ě_��w�o���$/��׳/�׾\�`T��U��:�|��Ƭ�w��͒��+�$N� ��j�<B��)/����j�r�<jl�Y������@�i*�~��b<{��F��:
x+B�c�f~e�3b�T+F�RHĔ*����*y�������\�k�d��#����P���m��Ei
�m�	�U�7��Q�ۚ]'U�b�μ�Bpd��/�"|I�la�)A�)4�9@��H�^E���@dk���kbky��*-��~���Ȥ82>%�u*�ٹyxVQv���!��<����3�]��EY��o�����/cez,97|OEԄ�u.1��>��;ƞ~�Q���]�5�>�H��:�F��P�S	���d�[]đI��.l�����s"kyac��q%�A.�g3��	�g'�0�� ��sٝl�[.�����\̥|���P�*��i�Rm'$>��՛-��we2|�Y*-�Cݶȧ���=�Z�	��꩒��4��/S&B� ns͒�W�3)|=|�Q�-��<NRjo`�2�����G�dv4�X�G(�#,��<�"�Ȩ�ijڗ��%��z���?ײ���*�.�bo|��gLj�[��~-�^|�N&�]���6�BR�rP؆��~�'�pY����c	cLVx� P�ȹ�Qn���`c�¨�Z�����Ϭ�K׭0�z�NF�ZZw�ΨmP���N�q�=�%<4�U�$�\��u�+7G�;Eڍ��[��Z�&�A�FIV1`b�;�PX���(�`^O��&��2X{n{j`��8=�qٵ����y��3����{[�JYL��c����Q�p�<�.��~�b�˴�TZ�F5���5^���%|�NbUՎlG�W	���:�/�(���ѝ��=�v�4Я)8ɯ��2/��sY�%��_����C��"R�[b=�W�?Se��:�W���acMayRH9b���DcIu����V"��A�Bm 4FY��mgZ�?��g�F�ڱaӣ�sF��i2̍��k����b��Pc�$�֑������U���*�Io\5��]w�![Y�Łs��uI��1ɋ�:x��z"�)���r��v]����L0�:>:~sE�{�ܚ�k�I�<o�g�B>~��Y�U���e`�D{T�ҕpp��j�cOH�8�uG�Xe�x���٭��q@�nJ�WV��NG�{.�ׁ}[�"M����+��qYL��7�^7dX]G?���;��I&�jP��kSN[����݅_W�Ě ��(I$��6��������~bhJ��4�����D�|�����^w��ZY'�7����Z�Y���B��KQۨ<������n��"N�1�`g�rs#\����ܾG<@(�Ϲ-���$������Y#I��5�$��}�ئc;b��
��Ԛ
�ZW1��;�i{��沬1_���i�39�;�F@�%]N�q)"�)���peS[��m^Zt�&�g�����aӓ(C>u�<8'������b2M���`
���2���?��=L�̒k�)�q*������&[O.Y������e�4)0��f�W��kx�L�??�U�O��UЮ2�Ԉ��c^�}m�怱pfs�*q���}"�Ғ���5J$C9�H� �w��y�A�S�U�4VD��K��i\�t)gRK����F7T��~O�=F
�N�BS^��2J�NP�x\Ή:��)��X�q��bԗ�w,QuI�ʐ���t��!���"��^ǢD������	��Gs���,�(2��̃�*o�fL�$4�s��NҴ{/uX��'74:�Q�Tx+��ԍRjM�	g����{14��`����u1>��c&��LoQ�c*����vm{�����YR��e�2N���4.��yI�s�w�9�\�{�!&4�r�]G4�m�O��ΎӚ1�`�/v�X�\��[��X��9��]n�ߦ�y@��G�밸��uVt���M�Q��y��"�{�yBr�2>���Ҧ>�:
�gQe��BZ�/��,a�+�Ln;�kXL�Y�I��4Ld��	=4!�؝��+ꊱ,��=��_�k�J�.[^��<��̂)�������qD������
�Y=I���%*��zO 1''.�G��8�GCG�D�t�-[�=d���`9�~����G��ɬhr�~�d!{�!�C���9o)]�8~8-�.�����fOأ}���Z/�yE���v�m?,��2�j�.h�i#���NJ��k���u�p��F�-K�ow�brԅu�������Y��{��Ifu�DU:m\�r\�E̮�JNTl]k�(��v�c�� �F��\�*�L���q�pS��v^:��+iY�-����CR���N�8cjH����^Q$�+{yV��m�����9W�]s���P;%@4 �J_H/�\�����4�������	,�l��0t�=LP9��,r�=�J�$^�&�J��H#�0�X�+�trYB>��]��e�9q�oJ�I(Mjԛ�����)���<d��_>޲�v� wV����x'D�ݙ|�z�dg��ݪ��O| �{S�oHd����2���Os�*!M������&������ �nj��F.�Id�PA����Šj�k����u�kC'�FJ��,,�'`��S�(d�b�
,�l]yDR[c��⤺�)oI��1�7/F�\���  ��*$�����u���S�d˰��'�i��:,��	�7")�,�=��E&W��:��+���Ǖ�S��q��z�7,��^�tp2�w�:�D���_��X�h�E��M��>���D�
/��@*/+���=����R�r|r��' jiC�|WP��Ɔ�ML*�̆{�g(f?j������.(:sH�W��[Y��,<���E} $�gc<�Yޝ��RRN V��N�ld _S�Qd�<
 :�D���v�:�"�?e7S��vo�-$�0k��A�ƠE���<D�e9�K=�d��7�R�@0?��6�?�{����!�E\�X�1İ�-�46�:B�I�د����B��n��\z������q�K�!B�j'2^Ai61ث������7�<!�7�{W"q	oUt��!F��յ��iQ�B����h���i^.��d1�դ�,-O��_�;EҮ�L;�E�3���͕@;���Vq�ズj�T��h���x�$q�Y�y�U��xµt�{���Uhz)��F�^`Ϗj�4K8y%[����}��8�X������t�b����PA���H&D%�cu/q���0Rh`�A���A�:�Z���V$S٭Q��?*Lx�N�#'��(���ˢ �eN��H��V��N�r=A���~�i�-F�J(�-���.`���<��CN�L�p�:������L�.oJ�� 6�61i�UvR��$q3X�sub�`QCʳ�s����$\2tp��㫻/���ì|�r��]���og�\��(�F��@���U��k� �h^��=������`iz!���D�on����U��T��}��a��(	���P�`�2R�j���-�O�-��J�:�w�w���5�Y�����T�73�������?TYbh�I5��~��A/u=�Eˆ�=�+�`d�\�4qu��,%�l!��%�{
�	w�y�
wG�����k,�G!�x���ٵ|�GKsvc>�W����Êĭ��Y��*�8[y+�$��|�,�$sV�"��76a|��8���D1
 UT<k
(!��U�u�ʿW��7JĘ�O���_�́1�$����U7jr����~��/��],��Fy��7�S�hz�w !\{c�Uvv�-��M����HQ���͖�b�l������MI0Н�G�z��>�	�G�>�>��5v
�`7S-N�4.�ivw�B�2��T�'��p���%Ikt8�Ư �1^cѤYR�_2�nV\:627ƻZ������V���ͲU�t����O�i�|�#ܛ�Z-�mݴ5h�Ĳq���+ZhRQ���`���>*�~�9e 1\��F�2Fx�g�?��6�#=	��=1�;�7����RP����t��y��^�,����DM�DVbPPW�Y��<�h��+xO�(�c�r��8��r||" �-�ێ٥<�rk�G��z�o���ƚ�P^�yQ��C��ߘU��7��tQu<F��h>9M��#�i��D���f�*|��X�os�Wd��	%�N�2�}~�hM�}��>��������~�ű��`G�O�\/%rB`
� "󧬫\ �?���u��L�V�oy�'ܽ��}մ�Л����/��xo��H�-&zg~����2l�
*�<d��2�;䮵B4�9�&�@���r#���Rot��R�߹ߥ�#��K�w9�
�_lVnw�����(9Gaz-��¬%nӭ���&����ǣa����m��K%"1�:ŧ���o"hn����4��e���:+�"��O��'w�B��呶��RV8�o$R숃�8\_�t̏7T]�j�	V��r笳�L�[",�1��MX��ٛ"GtF`���ő_W4����;�2dC����%������NI|2�G�y(��=� w�@��kv9c��"9_�d��g�N�<%�[�N�|���È�����6~\�@&p�n&UI�hT,��Ê������Kp��֟�\cr[�R�%�,;H�����x��@�9�"(Q	�-8�T|����4��/ئ�p˿�����=�"_�{�McA�r#�c�.�GS��k�&�PY �{Y�ҡ�$
L�q"%?^#W�\��>vdk>`@�C��4���]q�qvyʜ:@�����J��h�౲����GSU4d��X0Իޘ.���Udw�@��=��{�aD�ک[�a�Q?ni���j�bOǈ�����/��E����X&�mN�"�Ɠ�)���)���g�Ǜ�6�(HGs�,W�	vT}�]���x[3�_����NW(��c[�]�7�(^��Σ�v��T�N���o��r�T��?C�<��	��%�>XHi�=ö�?h�'8�&LKKW��F�t�	��K>��= �*�2��M��d��о�*'_��J�9�b�{u�T��,�u0�#:@5JdS��.-t�9 Ũ��F_f���==c=�tm���11z.zqM�V*��ca�;o	Gf};�MUl�b�[i���'D!e�И�m3��Mj���
<gQ]Ձ`0��}`��V�ވ��ϑZR�8�K����н�8�H��S�ג^�m�i��]]�<�qKL�o��r	�E0}؎�ϰ���*�������hF�_Q}d (5z�T��VU��<�a����Ff��cJ�ц�K��E�6��s����*�Q�Ah�=ʚ:�K@��o*)���m� ��:��pLL��֔Z�ƭ�)�G���T��M�o���z?�X�<�=Wn�a�5n�R7�p��*���\}�S����ze!ث���[0�!?Gi=�ހU�Qa�|ƃΛK� ΁���D�FCd�,n����B�m�����5Ⱥ+��\a�w��ks��x܍'�:���{I&��������������<{����Hz`}��^L����L�Υ�2٧�>	����K��}��X�������]H���O��M��2g~���Rx��姿V���5?�\�T¼-��W�ź�.l�C���۵�|����r��Bȸ�L�o7@
1����7p��+�Q�T|�ҧ�x�N��T��Z�[nR���ų��[�^�������A{�|�<n
��@ZW������yN ��tB��(GΕ�Uh�Bک+�)�?�X�~���%�)��z�%�b������/����s���j�вC�6D?�q��:�i� Q���O�h$��+����'�CnS�{q٥t�uI7j[�N^��bb��En(�E4�e���®�`ڃj�c�tu�a��㧳uN����(i�}9��o���?po�����*�f� ��ܳt��*k��>sV�Q�di6�JG9}�Hk���1��V���s4�
J���~�5Q0��룭��1����:�R���2��R�9�R�1�����ݶ3$VЯ����w�XU � ;�bMɄ����n��).�'����h��y�����儯�T��=JR���3��'��kӲ}���%�	�5���/.]�o�2a�MN��ӳX��SKR�4V��hu�U�J�2�� 8Xy/�R�������Du��~-#?{�y7�X�V2ٮ�BJ��wQ�_UH��ܷfl noN�w�a>�ï9�6ޡ���=���_%я��ȼ��A��pY�_)��4��y5���TF�|�mh���`�"g�>ѦfB���z航�i��j�Y��rw�V�Rc��N���F1��ǍC�Z�/�r�0��#��J<���Ļ�}h�e�w��eb�z�'����L��!r*#��-[�s�Vؓݙ��psR����~N8�}�����B�ޮ�|
� t����X���A�3��h�z�)�t�����7��߮4h}h�26��)>���T��Y�9�����s^���W�;jp;؂H
0b�*q��)k�9c)k�Y-s���6�*)�(Z�
�����S��^Cj<�퓭�/���Q��եo�AԎ�y�"~WN��^��j�h�0fɍ�$��,�
=�K\k��=�]"��V��,{SE�(�h�L��r�n��t�f��f�R��"��=x�_�/ �"TP롽z a=�lѹ5��3�lJXS>�S�"`sn�r���(�f���mj������,Z�hA �_�g"�^> �Y�:��~)��^`5v��X�����hЬ�G������ |��s��Q6��!ݧ��8��}�u~��d�Z�d��"���S���ї�35sc�j�!�f"	4�R'�Aac1�V�>�l�/�睫[�X�����r(�����Fؙ��uDA���:�����Hj��3��z}S(JV	��`+�a���q��g\dk��7�s5@!+#�J"�}��10u�����x����1S䆵���L?�jjX	�+m�ȩD1�(B��_�T��FtT����/�
g(�Kژw�|щ}���:�\�Z.1��a|�0���f�Æ+�1�����5h��@b&�pQ�\5��6b�#%�1���#2:w��ۚ�,6X ���:!"F������@�;�[�T�q<<�a0��g�^5��c2
�h�j���{���K+<f  r��lc�g��,�W\����Q��y��<�� Ln�Vב�B�Z��*�9�0�h�|{\�H�K�z�jgX,g�ݹ��^�S�\��Jkj��xCk��9V�rF�i�A�#x�@'����~X����m�q����O�6%�l�^_�9����' v_�-45iZ��Gr:���W]]�7dp�M��~�C���S�^[-�j5�pY(@v��mT�=�?8�V͠��+lb]�@�1ƖYR��HR�����Σ�s=�LS����[r��<s"��1�N����,$ǋ��S����Z�-`����~(H�o�씊�+����%+d�l1o�]S;�3�1���p�����|T����L���f�yt�%r����`D�f����DfL�r(�{Kر�GgA��t�BtbЦ�سg:i ���$��~�sږ^N��ׇ�	d���z�@��'�׺M3������"�tx�S9+c�#@�	�]ӰV��e8̈́a��þ�����7Y_3�����*D�8qE����uJN)�7�'菞.�)�P��.H�jJR]��]�U&?j�6�4p鉮!�=���{��́�8<k	rC����g\k^.�����(���]�1ͯJ*I���rS@�P�3�����˞�/�?����?cZ�UHO
3�9���tjo���Ö$�!#W1yԒ�8�ۛ��չ9m�����%S�s�ލbn�'Fr�V���n�1"�\�2̥c^���Ȉ�P0��z8#�У�,F�'*ZA�jF���$L$I���&�C�{�F��W�v�2�y�w�rջ�q�>n�7�s�Y3�cR<�K�J��9d2PE�|c����,�ϣL��S��bf�vQ����S����x���h2�_�n��m�G��eH���1��H̵��c�_LT���JG�PO��G��7���6[>��r��ߴ��Qxy�Y<�:60X�Kn� ��G`��nG��ފ��p�yꡳH�U���d��Q���5�%�U3�Gc� {�揺@�hp=�{]��w�鲕I	y���-������Lh�]�P��ps/A���ZG�j�(dǣ}c{Z��#5�۠�?R��r�.�JJ�C�D,c���uc�̀��$�<"�h���z�D���q���v�1�~�J=�=#�������yӓ�6)�1������)t�d��Ά�`�]�}���l;��4��huʠ�����OWJ"V�[��lb: �-�v�.#��^����;V;��yIC��ر>�vsTq�
C{�:�,3��2��,��|Eg��O��^�AG�m}ɸ<����<�jz���.����*J�¨.唱��Z!vk���`�<_<!^�e��:�ΐ�5cg6���3�� 2�뤪�UZ�o�l��c�����^i`M.�Z�>ف)�({:���7)�D�|��F�L�_��Lji�r�Ů`�H�TȸLA�/��m�gY�8��Vr�LS�׃kY� 7j��t��Ċ=�w"�X�t?��#k�w��2P	���-J9���<��Jb�5�xG,��9B-#�a�y���g�]�HLȓ�AȦOwƠ|�,H� v��~wl�`���t��ݶluQr`�0]�gz:�������V�bt�Mn4('�o+�n�z4cb�m�dg�c��I���^������f~GO��� $�[�U����Gc�n �ua��^�`ʽ*j�qzC6���@��2+�J��D��yX�>Ե�WVO���>�x�.���ل��3d��"���S�!�h�%� ����z�(���t