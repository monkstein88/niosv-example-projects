// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
VRkg6523m7X0gyrO+sMo6CtiEvWSp8i5CtjHgRdIgnddNBduI5xmVM/DkK7QamcEjNkZo3JGD+uR
5oetOIJcBKQIbsw40eTmC2TGg6bY1HeeNTlMg9pHyPVMUuvYl/5TPNRloBoIUOdznxHy0VVa0OX2
9OK20fzRfqLFgxWPXvg8RjF2zQJg+V1zWu9tOWP444hrzJ4ckI3Tm2+zW3dZoKTK6OAhCs9CN4YG
M+0q8sZgnkRYnQiJjB7PbA0V1ZqO4KYRHBpaTid5jbErOSKr0DR25dHkwEUVpbuvMyrII8a+JGVH
t6jYOZI8MmTeA7Htxgar9qEj70YxeMM57/5dQw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10144)
SwNaKUP3WrnlizcsdtJbon+ihxtTbbRFzq84BnN+sdseEBk2RlXMeuPHzO00Xx9OZM/b3uyoVIBM
noMiBW83+PU04bd9jx+jMNqwM0Nu6hiMmQauY3VbL9yTXJatR6NbK/nYnqKtFZxIrEPIyr8lIXAC
tkMOg/2gn2CIuC0Gfuoh4Ri9d+QzjkBrFSWdVWAQJ+xaaHuZ81i610ACQzZ5JZ36HepLIsPo3h+H
+zWltMCVnSMSUTODm8ArUZ9rz5oii28Prar7biPkHLTkoqDReq4PC2dTTDxeX9u2r+tPTTg0M1pd
eqQipDy85wdpq4dHizRVJ5Kgz6Wq5UWJt3oQTAx6CxeO7kHN9Cl6Z+1T2CVSPHwYi5MVJY0x9PRo
r5hjeDqFh4sGF4qCg7Kp0zR61FVcnG8a3DsaBOOurndWKe+a/0j8TSC0Sf0GokZqgBdKoQplcubg
vUt1q1p7zlljjfpwr2W04taCQ/FatExUDuk/6DXZXJB3axzABvlD868iKErHx93hU7zPVBh9OvTR
cfmbD5uUGkIcHCUHxJjZXxGT7ty4Wl8wZVV61h6wlcqOKZ7UqaiyZNNY6VYiYAwaor5fAHlDlPKd
6lgqRiD12xuZQxAa5mgfEhv1KVtxw8kClfPlPiwInfilxwZgyhd8yBuitxAWGz3KymVNgdwB8b5W
YoxlwkQxdYZQxIFhjlNVxdQVqaMro3kDOpC072Q5k4TkMWlM1bWpPT0fJYsIxIteKa1eiHF5Wbk4
cPfiVcS9o6eOHoyjhEqp4Yqe58Rg4K/6w3wx8JAqMPlO9uOjVF5mc08ueGXRO2kUnHLzgTGvUGhs
t+M5GJ96EsYLflV63GQTY0vSod4ix9ZTmycWQCM8BpnBxrVt1fvnbt3UveOIoZZvu4dgvgfJmpND
5QTJSR69BWjd9QhMlGzae3mpyoYvTMMrRWkCIwJKvKizwQctj+/zjVpG1YaTIVD6z5mjDmd9GHPo
tLzYevv+FnKP6N4Pfx2TmZgChr+dwYFCg6f3x6JWzR3FoCWiNFewxJ+c0dWeRXtEV/nQ0GYZw4Lq
XnbRjvn8RlOKnTLg5m2POUpk2WHdqWNK+Ik4AVqMevkc72xnsEDvqYqq8ly5bU5rIChDcqcCPOi1
YTZnUkm+QesHtHDJezvg7Bjto1fb9QT50zy8wzzN4iOyl84+FC7CM8m7LU2e6B40qTAun15H2r4P
2wb6KY7tL1L78XhB2ZqXFImcHXhL1uhtkp5Mgi7+TDNQmEQGlugKRAe3vdwJpwNG0VSk5ss3la+t
/mlIzvRPflQ3ox5zUkzbMRpiILZZkp8wwKc0OkAREFeMoXMc15hakv69W4MOaViK7msFjkpqSCLh
NOe+AmcUf81P+49cyLUM/eem0kSsx6N4ccGmr9KIhAi7jPIJ7QdfnYwXsZVvFdXKyaqWYntmkL+s
YelthSTYUGQ1oPVv+1jhfvmjvWh0ZKvkHnapmM7FIirqIdz0tfzOgVx5d3tXBuui15Iq7UgjT+Fs
vza/2SGWV+WhYm1RLamyPul5MCXMar1zUXallB5slSdvAa0QdGl615+LrRo+NVqWIolJCUUy6Y4M
Vsuh7ZvpwHt63spMXYbA/hG6w+kXAu+KqKCA+dOr3m3rIonmfDPa7bQr2hpi6Vur+vZd+k1jsgM7
vCDjYBUpZO7YXJEqYdZ36WlplJDaPfcwGvesx4/9sbjULuOJDTfuvUXQgOd6FvzHH5Fb6O8Zkb3d
FYRmeSHES+QTx46WhTHuAU0gEVCtudSoE+GfFh68F9pr5Ft9qg/3jfnnRiAxOHsWTTpNGFcDDc2Q
3TLQ/nyI8I67BUjo076erKD9UiZkpAhx9mSxLTjnU5k9v8dsETl7iFk2UMJH/R2Lk0hw44ovFeoc
FsxYkfJduywIWv3unojHatpxvfUGeFaFiRYS4t/gXxd7lCUzv0THrN848gdTdtfWH7iNytdDvNJW
QSIAhAZyl1hTgiL+JDp8peNkZ/7lPo315JqTXq9QRbLJBZbz6f0SppDcZL1yI4UzpAZtRGiO64Am
maxwBWiBP6OrCW7M5GsqCOqLr7w1+ZhPg9oTlmyYFaNK9EIVDOQ9l5AubVCzNZG80IdA6lAZjVJL
l4Iubmu2ZiAZeF6BxglS36IJ6QBeONbtkD40Iib12pK1V5I3hdq0ABET8h/2FqU4yleTVCSJ6YjU
gNwWLNST/4zZfkYyrkV/IHVnASzVREgAhvG9/ks0hLT71KE6MY6cS3NrMUBrCNvgY7FiM8C1nRsn
EYrxQbQ+EWYoqgY4hl/Rutgj0ep0u91Ao7muTsA/UbBNc1tzigCBKu2j2hmquA9Qr4bEZ0o3s0Fd
LMFn612Amqa7+bYELvfGYtj/oviQ//4ZpxUrCwoTzDkaCWh9e/8wDPJPLiz3WEy6YXYhFG6ppT1m
HVfSNJBVzfEOc4bz+0tlXSqzcaUHiI+BfrErbNMX3+VTKcsdEOJisBU9KCK6Xquod3HPdtesj/CF
NOG728H11+Ya+71Bs7AMTWE7ev3+UUVzXyJnRRc3EIOjBx8ApQo2ReaAE2zVGOXyBeygnZQ9DP4I
69aCJCvJF+z3gn/dgpttZsvv5uUv7lPl/cnpkQHGYJzmyVTHLG2pyhjROGMnZbuAH9oVpb4ZxOCU
TAD1CE1lMMY3o/ictj7gAhAPQWqCJgywSwbUmlxa04Op0x3NqGutnjiejswLaGt9TfjzCwYeMYYP
b9uv1czJzKEI/HQPqQbI13vQDTAB4xqPRdP0m6jztuw8zLyPOlV+Zag1P8mI+29W4bMdnzVBgJjs
M82fbleF3Yi5UqJ9sFZzTK410iP5MKuGdwoVfPldaREyrXsvHbrHgnNrGcx7lFnCZ50ViW4Oqhvw
hdccjt1ZUrKqMOK1aIP9oqA47O/ZTk0k67JuEtSAnFMwEPCWsFzXOqlsb9zpF4u1PxwrcHIm7opP
+/tqBv8pv5z2GGCCs7svJ/gnOwPweWrMQ0HD1uNxU2mnAUvJZ/CIzu1DAo5w/PMwJDt5kwbOMgEi
ulc0M22yx5H3eenjSjzlETdKpMzCvTV85iejxVar89G5HuRZpN8VDv0xrhRnuCvrQgSGRGDCywkW
GIcGQ3PBEJkoO+AwgAqrL5FdoFQEtUJEdfg3IXb9RRn4PWbMv8Ir1pnpEyoBVT3SjhaD9Wx2lmFt
FUTS0IFH6j3oJcwgu7cPTq3iVO03dhTKjv/9lJwd5r66ITxcd5CMjAqizNq9sW53lCZt6IVb7zfH
iio52lbE73WaOPtl5fGasPpHGjeutZdUejNQbJk3oZC7S7xo7TxDd17N2gLdfn6iPnj7YG7lhYXP
5fvPe61hvmnhpYJ1+Lwq0zk1Sd/yq2ckjcp2AETx9RCqwBrOjRDeT5PGIcjwfjqEmFLZyDkPtQSu
sJ+vT0KfGkSTsZyTKtuZ4Eh0n0qHnFZbyw0tr53iDzdBLkAdBoWGnN33Kq/FFIz64o8/1/FZ+yvQ
tORpHWNWJwX/2lm5dfpLegZWtb3WYfB+5y24lGfHUWIO1VbPsmG+bmUyBacwL3V3S/5gD+E+rS5Q
79pMNqJ3fNh3z5SjXxyZCeTtNdtEx7jDq9E4yzQhDGvos/JKVn0g7QWQtPnBA/f7oRtBAT094hpi
VpIMQ9yZEBTRCLDD/fgBtKyjn/7EobKRJsGtP6R7zZUdqfS6Y2SXlJ/xDIPahvSffV5K0cckPjxt
HQROS+aJwzudyX1b7CvhXpY+YYg0nHamOszNxcjc/NlXvpX2gwfUvW4bTkOV3zyDtSMHbl7SuPD4
RJtLCip6myudLdC0NYDwcHsn4f1cuszjShTCTKD3A5zHXlHxPiiRYVazgpEyjUib6KF9qW2gEARu
kz7Xg5LRwurxrnY7MenvzgJqeZ1RHsHxh2/0mlStBsON2jjjzu1N4pivb8LNqgd0UEBTtlN2YJ2n
vu9BsH9I6dnLMA5x7pNHDipWxEQha5h8aT4Jn3XJOoQ3imGNQv4+nG6s5udpXdAb8IhaKr6LJTaC
PeABlLlCofOnx1h2nKMVqwSqwcLl7qp6Gwtii2twf8xX60TU0la0nODi0zxrIse/+Sj1HylmXKOp
eWPmh1I8NoSlshKFCqjOUBbtlB/y26WnxEUJ8AzM2mml8Xanz90vYyGqMmVbp3Jbe2jbNGoC19LH
w4n8f8j6Jsi1f1oiyN6Q7P0ta5dIjesFvWHzkdRm1wI+wUCZu35fvuEatYQ6zqiFrk+GddESHkz/
PY+YP1TpSTtCzhKu/nfOcPK1IyC47ip42RogZlYHbw7MFMfrSu1e8DrHBd8+UorJHccEOdhvfEod
sv9wrsM5fk9JijLdRhjIMMrNybZKaJijM1IuQyJvblG6AmzbFqHT30Qe2SA75xsRiYLU2OwsgH/3
MWQUTDA5ElReOd1lGsDGqkLJdGEd2J6iqMPS8MZUXx63ttF/9yPeABpOAyKMKgsLueszvjZSgRTY
utVc1dHCf88icvEYidEA7g0Zji/VcbqJ55WdGiuZIyNrlJzVBvuhRXgJCdAYbIZSp4xLQKZbr1C2
/e0sm65SFdZsASJz/xPg5hP9v4IITuR5ikmcfbrwKLZrJ080eBgNjnQMZaO/fCjjB9nUYnxf0PcO
iIAgiSh26HvUdMbnFvTptbQ/x96IkdPorVVzlZ8zDeO6O8exldFgEFNaajQqaDBsnMr+Y3p+r6dd
9SP07wTMvVpcq+0/qhY+/n4/0RdaUvFOA+94E2TwpTJUw1sfpXXsH7Q6c6CXSKm+VSjBvfJYYyPR
+6sHriVwKnbgjyDkpEKfyDULUPMByKv3uk/HxCMGFZL8fSXOQ9Kp5oCjtAeXMcUt1MrlegPtQFkP
tONg/1AWKWyvOkL0nBlHE7XB/dR1bwbkyyTdgQTusxvz5oemr53+fXEATERil44okK9obrFVPhkl
xTXqqX3P7xyhMRVhkAmAd7u59mTUXi8HmHEFyjUNvlz5Cwc69LyGW/KY42ZtRDLZTO19Utkg6bMr
D/JIJV+NCo/TPmzEXa/welgk3yuBNYXmC9JxgoQLJAPJqzmugpJ0p585xo/hELMdN0FSg7xt2bxD
tmZmO76xhNk/bab8bLD+SZI2SsR9n4xncW7H+aj1FtY8X/ZKIsFWVkJj3+sFSgkBZfVZnvopwLuk
9cxwxRH9JVsJmf40/c7nGqmy65H78S7++kC2+xb7dqlKAcP1ctbZyH4ngoNFT2cpuMivuygtO8uM
CUn0T1xTihY2OYowNY1ZXuGbWa+b4/ygVqDalsk+ibMQxdRRj37Takp+PcdrCn6twF07ueLhWQSc
hFcfO5zQwgAfFU295JxaYNt3G3s8AQKiaJCouZRdz9gCB8/t1kmLC7P4YbEU7I6mrQ8utKHKjLY/
BqcUC2Fj0WrIaNBC5YMwXuj/CZpeUixKQ9VUhOOHRXjxIwJ4FFedN+v0xtZ66qh1j57XzQRf+R3X
QLsJuuOo/zFpDaElWgpAX8buE51945lYTl9Qrm3sKfI2qn5N0mscMnmYV4vNWqnRtC23o0jWSbq8
1tU4TUDhWeALa5WW/wm90pv+/C/CacX9PCUlCv5M7OjP3ZXdI0ANoWYbSvm56yTGdyEim9t77RLo
VYmKPdJC+WaAjQNSv6VFh1HNgJLmp+co78BIMuQiNILzK0x7YnJDDqOGEq5IorGaO4x1WQrJFDc3
1ydCtB3xj4471gEDpQBLQisICD92lGKsMMAapzOGTkpTEKAZb5R78j2liJtUzX/2Yf9/elD1VPEj
CPYiANTS6GOCes5txlT601pGx3XPG4pL0NJYGoc2lviDW2eoqanaKPZRN6R7VE8tVmyLy3SLkejS
VtJ8jO2fHYjHoclT3A+D1TGD8xAFhXGr+93CmAUmeoro6Q7FBR71PkG+06NJVPMNJWd1m+Wl943E
1reSaMmtBbtb8CbF7DtJKhG3CxDmJeKgo8bHDqeofTncH6cM72qhsog9mvMYILKSrLSu3kLRtblS
O1P36FsxHZfrQUL9YBgU9Kp5gfHXF4Qk7xNbr0sWPfmdBTv3iZWmjoOdI7CYQV7eKKPd2txcixek
ZX/AqMMcDGkuFHPYAB+onIYqjjTKrg6R/GtKauvr0KETHzXG8IekUDxhWs8qQO4N/IOzcQ24vwmi
OuHmhzuMCxZiD9a53IB1yUM5KDCVrDQsmav6zCFGHk39tSIIjBmIuNhh8sMIbN4buEvgQGBLstvL
VNIDh6M3+bOO+GE5/fvz5mYrqHKlHMnEEC4fyFIUbqZX2OOeyq/Kaa0kKJYFahqbxe7Lj9EFepdj
6MWusSkA5+/kNHJHOZYeXNTek3T0sqALCZWd0akHmHIuYwgyP4vJW7RA+ouGSmGeZoUPePhNoa5E
0XBqpPDKNgNo13Y7WJ8JXxnPE+/vKMkwx3Gmr6XSDBacmSgZbms8tzS6kYlM12nvJrNeQBQHQCqm
dTmUJ0lbNjf5h3/UUeA8kPWEMbr/2tiCKYoW1BWlIUMBW+9fqnanHTYmjmfdSvhj2NOtH5Da7CrT
7vLNsECRjvv8v67oFBo+UX3PtaLPV5thiyaXdc480fNc3DUr2mnbI1Wx73Uv2UUETBnGPGPFTe4U
P7uiTeLvMndfjWzqwI8FBE8sqUyOG7HvBhvyh1kTOQhimK8hulQYv5NX7TLfqq9IKduMAGo6PH8D
ymQ3zQU0y4T1W3XudXAbX+svYFoYPOfYFmrRNBnGqMwPtG9imBEmR8WyVU/xwkVT6VYWBZR5p/hi
SY5xBQzPVmpS1K8YpfkaiEK5tvbfvTm7KQ2FE44lA+p8IeyWV7LD9nWIfhAVHD8AmQpOm7p6bUt9
CKT1cPPQBlJ+XOdel4JqHLXdISSmZSrBm+gSLY4kMbwk/aMiPpmgB+SegVApif2mRZ9CI0G0MxXT
X0uq6uIje2NQqM8TcLYRi42ZDkGRKqRX7VuDXQ99YXG+9si++sUooJEMT+yLBGISYlH58rwQXhwa
pmQ2ae5VL/+Oy0ACX2Gi1x9H+Zxfz5D5y2KfyLICVwpBUIWN6974+NbyuBvEGM8MWzPUotoCC2LA
NTCh/SRf5qLDaea2ypbgaFMT3SOAQY2Uba6ZoycsbA0GOy9VntAwgz8sZeuvvlxBqCZg+bYDk/oW
VftPGPhOmDnPaeRn303FZ/5qJPbx9uCilu8JBxNX4wg8UZNhTRgUMiAkgCfXlTCSuMvueZpNzBLq
RAQfJZHXK9GacfKmyYcMCXGMdokHQO5LWUIC2hrp2EUZXE/FNAmBYgBJ9C3U0PoYxRYdqjcNccsX
cajw76febicq+2CTwRXzC6g8wNqx1sFtdcBcNb4CbETBvkMruSjZQ2kI2ISJ+mrp1UJze1vnlH5M
d2POYUXsQ+pnrHeg0NlyXIoGNhSjyU3Rt1egWq3eU4i+vrSfkT1X13QGTxuB4AXptq1ZsW4/U1YE
kcyxrAxtx6CJ/SjNDjWmm74axFcLQ8DnhXNWZnSv8kqH0Y+Uo8+5ZJo2N1DXIU7oFxDwisLO0atz
zo7SkCmwUk3DY1MH6Oz+OpXRMyupEswUl9FYSX81Df+IQk6aQ74oDYD7uV3LxDUtGXuQi572GvCx
6nUWuLYsFMOHI8hG40ACSwyKxrEWC0FQ6Bol2idFOh2jAbyd8UaRnt+tswJxET5pZEnmyrsP0c0a
t+sTTO0G+R4e5Uqc6AR6tnvGb7cYwNQ8ScEuwMI/huKh5t+z7jW6VjDt5tINnwRYEphpm4QpCmP7
N0rqOSWubwHUpSZXZTPyd77HBcPhRovRHNXD7M78hKCCTl3m4lcY+TysexKE5CtCURg1hIdK4YT3
bQt4a4zjDU8mKO5q+AmiKUfYPUJj/u2pprzVkAQ+xWvPbhbGek2AYLSszU0WJkUdnRPCaNjwtVus
QGbJ0CdbZiWU562uaGUjcYYBJ6Uz12/Pca9ld+0Ij9oTUct+n+1+Xts8dm0Ajjvp64BMmaNVoRvL
xjyFGohU0mmKaNcfS/nVUfOMZMFt6ag2/RlUVRmWR/FA1t3wwQ5UsNjtE/GmHxXh3Rhdjs7CyWb+
jkhmZ3m1q70ShhiMAsTm5mzytpozN40SS2DU9sqdWo2zOdbMoB21VD2ekyct4dnbwfgr9/ecDWX2
LNekiBZpb8iuK902zEKLG8QrAlfPo4kLdOY6ZHcTCTib9IhtTy6QwufEN39U+FPDiK8MTsloJjqp
2ODWKOF7ulAZaifLmVAKmcWI9T1zghakdjF2S2zFHUlzJDpVRzKl5YZjPeDZhsa6IL3MGoQ25nZk
SNvJ1sctvDdsphrzPD++p/kwi7bFQSg3bfKzI0Hys9v+IPYX+vcG/YglT8lsbOAAov+31tiZFhmU
QTVwToLpeqNhmNj4dn/VXJFWvJWD7QDzO9Z7W/m5AwpIv9avAbfK3ZgHyOSDaiweVAJBXK/p8eGT
VUWmf722hIP2/YArvjJN0m4LbvW8vcRANDtNp491afTdOF5QFMLKg8wGplGRErGu4TeBjfC3MPZg
4oly8BrGgJXYBlR8igs1G1F8qbqUt92irafrJgDfJAEYsOw2g+k4iyM/ujatdX+P5W73+fK17IIW
3TZpWy+3gxbUIF+9VqKlvsBuP9FNNdK69H4nJlYLJGSvg29XhUmStt+3mJs00oKusb1HGw4E+O1t
p4Q9Vy7FXaavZHb/sb5np0I22maC5BimQyfh+0MY0GfbiKr/AV9yxSUZsv2QZY2jxLLenYAT3XOY
D8pGMUpxG2OWRMJW5pqtB/PmXlE8TYytJp4yj1CGf3q8wYPvkJzqYCzOBHkHXu8yKQdXlLTntV5x
yUYWCMygmSdwMG7qocwlguGF6dFZqgrO9X7W/M48A+rtbsKf2xoD472S6NzE51m+v0xkGfqti1XU
bbhvQQBY73UT7u/eKPTnNUiHIJKedF832cInsbxPN4cwacdGp+lEwFJAYbbN0MaghxQ07DMgRy5b
Vb12vLSS3bDWG67xBHOIKX+dOmppZGc1l02cr0mR+iEJq9yugQe5soFkwqMpRmCCsxek3297vSZn
/SH6Ier0TvGhQz+ZRpPkIdOQpfGB7saNH4jf0DTDtvji0HbSipo5kyygG/p1/UTlQsd+vZbwkNOi
ITQBrkA/HJKulCuQ+rxRJ93HBy7al8tfGRqc4LXzX+4tVrWuzu6KHE7ci/d0PkaMu589WkY4+2lY
FivwlXy5ceuleFr7+VL5aZ6MNXUBWHye0zV1+viJI/BSFz71NuDRo5OIdqsgWZfqxoRz1lz4HcQm
qMXBpE54j3fToQhBK7sqJh/irC8imEt2VBg79dHVxYmQmt7/81rsWdFKn1R9IIOLnTCepjAub8sc
HLPSRH2CR6es+OhCBw04dJ48xAPpSyQiKR/07bz7A9txyKf3Pv8lJtAq6ciW+v39Selgl+trZXrk
Qkn5LaYb5N/rAk3rsjzK2o8+IcMVoPOwNrQYTW954FPn1jUPUVxVRni/8yAKpM9X/8thG9zo+OPM
ebZUrKrrDfSaAL4HuZLP5F+9jYsqLeCtjjQLvL7l6ScYw30CzYPGMbbmAx06WIXpwraXD7gfYOWs
Yl/cMT0Bf43rjpLmqPx2P9ITLO/uCRgONPPqlQXM970cZ6C1aNq74s3WpzLndJ4PfWeQAfVs/mzY
NTBKLm++HXidZu07G4YaNDmjdNU8deU4laONqh1fPqEb8pD9uRSePhw/6PRCZE3c9SswZ1hawBKC
3ZgQ4v3myej041ecyXXV439MtSPIiaPqVZohUhNposfWBwqbfRUYSEXIh27nNC+8ccgDwItMR7+w
jkmnDr4AyGMiM3FqK0Gc+DirqXood6gwI3twtEIobMph8HWY65tz+pjvZSU0OktwdDV629m8vMIy
0gG5ZCxjneT+jQ/jjd9OL7FtG3MtQ7oObxXgvYIPaLTcP3ZThdMdlx2jnt50UjQWL4q9Yu/4SyLH
HR1sltRVoXGIUkfrSsn1gubxjTUp65bPfy9Yz0uRwrvWHl7iSPFZfDFYo/bpo9M1kU65dDEnyspe
DmhLxi+g2vaahswbilze9BmheIZtjNPSXBJj+bcBIHYVyIsK5HS2rLY0tK/aFO2i306gJpN0Wmam
U1wpNpQ54ZyXxy2dvQpez43EAWgEq7JYg0u4VU3njWeRWvHgPL2jK1o8cQjePKx/xyzWNe0dim/y
nEur9VkFFtRfBJt5UD4Z+UYWgOQpPvGXPUsXu4h1g3nuk8DFCNg3dZd/Q9nGe8Ql78JOMS1ONOQZ
oV9Pg3Y2NFQhh1Bbl72uMulQaQqZc//G2imlVaa8wtG6tiB+SE/tA2TOi8471bfjCknfIf26flHP
zqsZqlv/wxli7sJ88hTiibXHs5q33cS+rhWF7lxV8gX4U3yBtaALjCcl6QJ0baPoFG74neBqSAez
3GQg5rdm8BDlj5y015CkfpAvW1eiV6IZ/i/SDmdOd8uGnyOc7ktEli4daVjqP1kJuQSI5ofqLCqK
U5RTqMIO/jML/deeX6eeEmNZvnnItGUsROll3UYwtdvEi1N2lcJkwoGYh24Vx8iCCMeYTaunhS8/
NEpiOec8hHVYXydBlKcNNzAv7NOQR8bc7ujkOFcCJEgmaBQa1jIT1w+wFiB9UHieeFUICxQ4znuN
i683PcR5rTwVmVQHTKWUljYoQOmVGPoShGu9zsXyFYLMJE8iIctMCspz4UyCHLtHF8j+FTiKd29J
ZP60obSCUAEEpSQ2KzLUKbux2FveH5jaL2TuI9DT3HdT5B9+ZmahAEhTjeHLXriaoA4xQ7jA2Ok/
SLej5maQrxcZPc4gqG1O+EHlviOYoyOTScISPS+MiMTBOjKa39nP0bnm+Sgq54yYMhyk99L2+oHx
4QfYsmwKTpv9Z5ydsJ17B2hZ4NAUwF6U79iD23EKO0d6ukTbsmSDEU38s0tbOCjltd6nmt9WHft4
9QwfM2gLwsm35WZqXO14qE7Drihr+98QJ14XvE0q7iBvXVHYd+HP6aL4xAqWiHOx26BH4ki7BWNG
lL9ncMX0zgkUtnsc/mIxlDRkLFE24BfURAvqG7r4PkwcU6XXkcPXtvreVRhroeG434+PajZCKjOD
ge4kGLRJFxyctyuzQ8rMnkMIhOU6cuXfcymVj2OgPmCPwzRhjTuAjOnVQhifxN2+xOlhMBHmcenS
QM+WHeuVPAfpBva+NwVUO6oj/hy5As1gd8Qxd/ekPnWSB5rjATrqoZ+2fjmkiShH3k3HvHu9rJC2
9w+c3S4Rcu/eckp3OMjLLH7vl1eHf9vOaoO962r1nN+SxdJmZtwEAuTK4JwdX7ujxhHeCMso3NKc
So9uR7Fza+3bQd3s/blJkBXJLMccAbuhKsK2qBKcwUl24qxKp5HF0/9qAF/OlBc5q7WWOoO9waDZ
wArLDa82PdDFba2uqUs4TmgeVPCysTWDMyzB1O1oVmfKqyyiwJJslR8tIK7GKI+1GALNTtwMFgAs
LAvBDmbyNRxdS3ns2F/WN8/yijLeanJsKDA4L64xpX+pA3QkQ4ubicpkwQQHf/Vgk0yqxhh99+Cl
d2FpptyTsEx7m3CjbwzOeH/9S8Ppd5XEbpx/xtTN3wPMPehobxcT9+bbE/UhEB96Rs/NL0+ARb4n
8ff5xMD0+bcRgR/Odhp/sb4x9XsojsRWDAZMf8+SwYwkjnMCMxlDgnG+O/NJqcwlE8vUimVbPqrb
gBl7PxlNig4ffxk+gWvg4ndsELGY34WhidlzouPEdZbsMCS9ICj2vXJETPfB8JFDjwqQoC+rK2lZ
Ze6sym5Y6Ie3/t+AoOfM7E6AwlXsteQPXKPjvlSNNV1AiitGMrFp3EWjQIVwxCCv62ncqPBjwF0+
G1NI0sFTGn8KEUMGyBtUSeQlzEvTTqB/f+m+WG14IXSjQGEq5mm5LSiMBAXS4xxue4nM77Hb4/nd
wlJARe59znHRFdAzmpx0tw33lJzwWMLvqTyoacPJerI47FSghzK5w7f//0vpivDSBMzas3VHXphF
UodKuOoOKqfMmMF2hiO66pRj50KrLI67F3YZqpa/Pm+A/BOB7sX6WUS84K9WneIuOojUDy765fB6
C8SSfFwzHaZZ4x2daXyjBOFBf6hcdnP2tfg1XSNtDTDfUdIXV6b6E0EtfyMfERh8A0vwP38adgsl
OdSUHmZDzEC36lT4Pr6Ps8AyZY8BuzMz02nPs+BTF8yIjRHc0+nr4DPQgKaVhMckwaTgZS4X+SMJ
3W8a92aNKFyIj/ATwr+3CkH61DxBXUh+6qLtOOTb/rTEi6fVX9C27E7XTvba3RugKID4WXid5M4N
R5teMxyLglx8FOt8cvSWzcDdExVzxlEsbfpi7Mm0ZBOI8/u8GmuA3xWeDkT+WVv7L64F6jWw4eb0
b/sr9tI++X+eidJ6gcui/YMSldviZGozN0nYx32/8xaxOQk8Qb0ZPz5aUAyAwlLytQkDDy3K6f//
pmTJCT2luHizTKca/Kx/1n6xKQrBdBINReufIgP0Zon/wCwgzJGSyfecLWdbTvjscqingdrb0SYb
s93/WqZJ75tPJUBPKh/tP7Em4SoHHedYKhB8uN1K6OQXPc0vosPOIDn41Mq0CB2SmGYW1ijBzi3a
KmnA92K4lct0tW7vzAuwoLzCREcCbnYz/NDwSqqFMGdZKLpDb4UbJGqVp40pbRi5QS7pXsdXO9WC
HqHfvK9DJDjpYMSdX99RZEA0roCX794g2voz7Xq2XyHPEakW7JUb14LDANRnenmQXhUG0b7WTEbl
QxxlIs7TkQ1EQkqTi7OPiBLeJY3pvwC6J3TdKRXpxlTNtbvok8aBo+vANCFHCu2PgVk1/gLs84no
/aCItVq2L+UktHL9Hofyy9wXoa+Go9b2KbNt39vIU1JE6RnLuPQAvZ09OlutRrLXbAeGFaPnB8+W
J82X3wBLITBkXHVEr5fMq4V7ZbanLGUjT2WjgbMQkmZM7JIwEs+lLsLnCi33leXuQW4WkoSz+ON/
L8hPwSidg/hvpt2TjpK9bYQxO76n/7n6TdWgFaec7Tb/vex3Pqf8IfnNMzQ7hG4wA62L6h91UNQ0
7xe5C2ROzX8qNBUxddT7UkQ07vG+wt5gArBRt9lvIXzQEz0X0VS/arGg0+7cL16tIPC6uhUXWlUN
Tg2QIjKlYcuzITIw+S298/8/JYo99ChLudzaE0Cw4DUSfLReuL4Wg5Xd8wezjszBlaC6yXj69V8L
zw4enO4kj3T8rpn1IVn0vwIRDc5KrUm/he5cTVAekyCiD0GP2EgVp7fWW+eRflA2+PDgQeN6kUPw
3/LEO7wC5ufawb8hmurMReerLr4SfIBidOmnAVlCOLzLRzrqbSkSQoxO97LSWc4xNccn82ktMpBS
NSKWEm85HJv+fIAiHlO+Xo4gxd3Xt2u80DJLAXK83SqUAEaT7xvNYk8cRZHePWecqG1FGJN9l90a
BmG2jXRLYzBf2zrg5nxUd8A9ct643X+jCl3TOlszKk8HUOVmiz8NZv13iBtK88F8R/2SRxV0Xg==
`pragma protect end_protected
