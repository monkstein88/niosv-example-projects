��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2i�>�|���B��,<��\ ��W�~��O�?��K��<$џ_�!�ʙ�EɊ����JtmW#�[��&	���O7���>�o@�K�oM3�-��š��Y4H����2���g��Q�<�[�rF�d`��V�)qǊ��͠!��U��e���V�j�i؜F��n{oW~������qUh(��S$�3��w������룖/�9hw{b[;�T��W����$���D�'���!�6�_�!N_�yk��N��Q�� }�ƚ�t��E��n���.䋤�ƿ޳���~�%��}�?G�]�~��fMӤ�:��y������(����.=����#bJ�+�bt?���g'J;Q�E|^^2�۷�9��,�-��\����2�^J�)���ޖ��ȣ�ϑ���΀��3��0�5��<�#e�([h�1֋+����6�Ax?�����9xF`	�N��)̞HO�(�����lMٜs&j	n8e%��Ѐ�&����|�r#Nj|'kkٽ���a����<=|c�m��;�&��Y(�� ��V�:@��I��F2�c���v���L�D�̈́M�P�>I4T����D�yH*T>(,��៪��r�g��2Б��qbU������n0]\�յ�a��Y$��;�M{�@Tl.$�^��	���>�� ���,�_�0�kp6"�������~�B�[O<i����m��^�Ѥ��?�E�ӊ�H����P�V)���	{!_2�mzك�����qH(s���5�����B��`�I��'4QS-��,o�"�D�(��'Hl���Jv����0�"��ЗiM)����qN\��0�2���В�w����!�J@��9=����E�^2�/��2H�/&D;"����\����	���]_�@����v��D6�$�"1�>�|��_�!�,D �3yhO}�_>S(�Ի��ll>j<h�d���K�Q���bݝ-��3���'�_9n���n�^�<�_�<�RLR���ܷ�t�tR�U���A��{�d������+��.%Ew�������$�,�랡��>թC�����{���b�w����Ѧx�B����>���p�6��!��D4��z����Y*�ߜ�揖A�g�{�M��ը� k��~Փ�\�Кl��G��D�Ʃ�T}p�T��X�sW�U�����}�[
:�^�������3�F� R�#"f�oiGM�o�q����s��O����gd�u���0���s�F�&+Dx$0\��kw:���(���(��p��� �Q�k%�Cf1�:|:�b��0_�X����aɗ q�"�#2RjE���1�!��_?,yVG�&�D�];?����Q�R��������M�)��pC�N��?;��a,K��_}/I�c����3�1fC��WҠ����ߤ��W������xȲ�ҧ�H�i`�>�R��4���)k��z��@-]����L�'�r�}��s����?h�{�4Ί��`z"[vψ���;�yZ�$�s.KM4��, r�֘��#������]�@��P�>�^�� :��ku�ڍ�-?bU<V(߭ �#&`��P��L2�X
{��dl<d1tTƗ��ᄀ�Ow��I�
��b�DP9��b�K�c#����@:0;��E����w��zP0��9#Hc1��<�X!���Vn�g��%ɢv]	��b��~r.G����R��n���^�5to`�u=��s���S:���P~���"�eS��c�|{4#$X�ps��R'ﰶ�I��S�O7�\�ic�u� S�p��p�T��NE�E!��Z�X���jR�N��	iXJ���3�[N����Z��<�^��q.�DY� ����������'����/WZ�&��<�����|�ۊX���caB��!ʒ����$�L,�$�+6q��F��/��1�z	�T%���Zf�jG�Uޘ�N���<xk�	D���8;X�K�7�Y\ք\�����Rv��p�x�b�������Q�džN���t ����JYd����S��]n{���&E]�J�:��qn7,|�]��%���Z�̝��A���ܨb8F6O��IK���u�:�hï*>��;h>�*\�.���?A�Yj���Rh���*h��EQ���O=H�#�L/�jS���L��������C���)�V�:�{!����cZغ� ݎ)[W0����Շ*4(�Z!�L_�%�cٻ
�
^�1d+���D��x��G46$����ꅨ��n�������e;ݽ</�+�g���G���M�T�vf�����T|��<tU�}L-{V����/���E��W�S�^�<�Q�=g]1�y��2�i�2Cf�(�룄R��&Y�s�s`�ʹ��b
c)����(L�ݽч�V�?:��Kbsٷ�a���+_�b9P�c�l�����@��ûl�è�*��'�|r�y��Y�N��o��o�)�P��_��s��l��
p�]X�BD=��2�X�6�I���X�� �Q��i��Զ;����K9���vb�w����-Z�vw���<�mϻ!3	�4O{���jP�ǚ�,q�h���(w���J��=%w���\��rm5Y�M��r�1��.w��ѫDE�}-.�"����}�.\�H�$��`�i	�����V����Ԁ�����ɻx���G��K0�{��~��$C��.V��%,��R�%r;���
�����T�ɦ��PPY�KX��#dO��Y*��^\4�/2����0K>��:��Qm�P�k��
��Wɏ�A�kL�a�CU<:1jo,l�ɩ_Z���j�/Ƚ������i5�t<d��W��2��)�V��� �*�WX��y�2�Lrn��a����.cs|�N�b?@ir+%��za)���/.9t�lO٘�q�( ێ8�*�� �ۖ�X=��?t�ە3~Z�%ͮ5�?��_�@�x}��?�M��#[5,�	�(*��^c")8��j��s ���=mD��Z3�9-�Ω54N�`b9Y��$�i�
Uu�0gf���&Z����)1D�|��~]`�.�Y\2��A^j�L��%rpv������Vl���ŋF� *ۖ���'��)���39"�b��P�d1U��r�H�����6�]W�L�H�Vc%�,��-�dWpe
��oP��E�U;�@ʮ,n�]�"�P���;f�
��`�][R��'��SQ5��Uݸ�
aϫ��&6C�[�.j�c������2C��à�����#a��m����-Xy���I���a�Gi�'T�"c�Y���X��^���X�6Dw��������1�S�C0)�~�<0��1��.��&�[r^��X��zX8��U�g�/��fq���e fq8�����)x59�K��ΣPXܘ.�����P�?]`+Y�VʖG�`�u�w���Jӵ\�Y-�[���[��
��>��ZR�FZ���� aE����� V6#��M3��h�3��f����#d��2�)-T#qZ �J���Z,��o�����?���anRSxSol;�0�i�AU򩌩�n�<_-��~G�g�"o�v��HA#f�n���mG����hτ]���<8!(]�\�_G��M��s�P��#H%	�`���(�$V:{(a�oп���X�[���_0x���$��9xt�"M��t�/IhiU�	�{'�lb,r�W�^���m��"@�V����ȀoQ���Y��?��s��#�\��������k��Ak�G���������X�So�k&��A�H�{�'6Ȯ.��CB��7e7��R˴�M�uK9+l����i��ư�3���;	�a�r�9�[\'�?�j�