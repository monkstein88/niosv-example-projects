// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
bAFm0Q9H43Srroc/t3BMkXKG7oIdkQnnWNnS6suBD6ExIV3pegzuG7yBRA0dPIrnzs56xtpbJUnV
xI+Bo0zxyVv3nDdeAFcGILNowK2mbj/jnpi5ZD/UnEkk03Bc24UP0iYxX1D01Ign8YQlzlZPNSPA
GzbOAGt5oCdIOtVU7aRb4FXDd5uLmsFqSGB+AEen71CRWhf/G7/Rxiw+L1xazfFaKqMB815cqdo4
TTddByN1goO13Z3zEuF2qKseSjsTz9L84gXb7AEYPJW/UifAoL+/LZXslgAlrC4nSs566XyZDkFf
AxPmQnCGJBCT0j4KeJQC8vxoAudqLSrP6HOYYA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 21360)
8PVEfpdwnxRDkAUgm47FpNpltzroDRNJIwmgVwz1ZufTs2kFFWy05n0DPd3AdF4kQ8tJIBZGyuLm
1p+WcAKetAiReCYM5uBZOTXaRA5n7BwG6WdONhjLYDXEY9HuYCRgYJFGVQtT2rSKRd9tUP92ZPKo
qRtix8JAA02xFq23r/Orkj61Kg0FkWDQoxh/M58E06iBWbWHynFamkNIgZyECuMTiqpqE2rwDUmH
ZoxOCmFtP7u8YKsHJwUiMPFyKp79OUu+6R6aimJnt28+I6fYT7VnGq21b2nQNfk0GlwHSKfiVSVt
OCksYNvxuJfAE4WvsmXxup24MCrt8kJt0P5mGb6KpP6iNKMClrg/e8me9EWTNeZtZkWjvK8eWS8u
5KcfrEJfjn+Epw7nV37+Bu83IjQf8jAcTQB9q2SWk0la90X8UelTlITZnYxmROuJHNi1TmVqJpQB
R7KK8tQGcLv8gJha/jNT9X/YHgNLKroHn7494R8Jpo+uMrzFlflGXYWYEIjtmoSqAhsyQUpey94t
G/KThd3ga45H3aQf+GAUdNEUH2XB10AV+RKxqhja4Tp4nYGeqM9dhUh/eog2z/79nHEj7R5GpOdG
lv3oe9ejep/Gwuek3y/YzZwGs2B0cobQzpNlM7fwyayMTHICHO/JhsPctPtbK9PNMNK7aEZ5VNs0
03EkHHF1DS11JI7gyO/X785oh92v8QjuDpvHfJqlPAZln6ZojZvczQVZNxdOwGayE/XzyN2QpxOI
tPsY7l7Lr2yBOBM3m7eHBwFNm273t3Z7zmGCrMtS8h7jm8SWZ+p6PjfrWesWwD8nTx+CKfQ26Bpr
aSsxa3wsEK2nSy3EEYa00MdaixrBoGFa9Ytm3X9B9Zho/GFONCY1anX0UfW5qftOegyjZEJx3TGx
P9EMKfU2IDRgXl+w3CY4HEA+9yDhbgbIvhanhzQWKRyHBCVtRz0T3+qY2pCzADacLllp/Px8UBJA
Xok3JLHjaCmpBN8+PPhJq2NSXkMJaN6OEXmxkaPVpnC0tj33wmWPcZa0fmy9iZD7l1saI/W82GTH
jnURvAcM6dgn3yy8fYcxBuzvvmDl4rLk9UTkTLLOTkCjEDySu/YZsR6wkE5NNWum1+bXT2E/BaGF
hR9zlq94BGdtW8hRbysSZSUIEAUV1qEv/FOCeSTzUnUNBWa5zroHmtoU/Q/0+WifgNUbZ25eI2dF
SB6VHakCox7uSVmCoV49esCUUVw4+4Fa1juQTe6AA/AHMamSIsURb/aM2o6wTSufglQ1jxFC7pCY
vKih3hHAxM8USLJIwmo5Y8BnZxmwFqJkjwejFUv0rcGzW+GUAyFOL6oQd+I/EiZ5XqmR7iSu1An/
q8jxXCxXkkJVBHk/8wsZc5lXruA075GY7bruP4AEFfc7K7VM/+KQsLhDTAnppve+CVDwNN2cRpXX
Wi3yl4EzWVjLC+YPhMkFcQi1I3JVHYWe6hLYFFFfU/dW+zXiC75VMAdMFWZEZV8qiPn7Wptw8WBz
L2bZQkMuEz3RO81sU+4FjYndsMJkmoXMBIJZMQ6DAkI9aI8B0h862rZaFT+DIzfS717QldeDktO9
CZDOwGtwbNazvvIZDUhHZE2mNC/XBZ98ens1UhRde/shSg0OiK5xDVRQQcJBK3ACwwUWXqSbcQrY
ujt5A2CU/00qFboDpsmm7if+i9CSQAtGUoqaCuvYwACWvBwWD7rHxwVPIrkTOlX0kGxdtqQYuSV4
jtatRT0BNR7UJn2FQ3pHOXTtwWo8N4Nu0zI6KHfsT2shMbCMQ0fcA+uycL+CruPunMND8FxdfqvL
cX7rUnbpQGwU3KxKo9PKLSyLnkDq4fGSYNr8kSZ0CaO8ifKHNKQ4j7VTYu7sMx4GWH4XjW4mOYrg
nddvqNFKj6HkYYz8gEEQOqZpDF6MnFnHG1Bzj2WUs2evFOg2pHKCPQTi5CljvTWQiptQ2VE5V+uH
njOYhlClk0lvR8lu3H969nPXJ2qrPZAg1NLtwVppjtl9/+l1K+uq7HS6rhJLW2VPKHSbFKXWsXrt
WrZodg8tN9XYBHpuskXetb3CCVGAA2JT2/OBm5gmzLFS0eyYmIIqlVwJt02X1P+IYaqnDcyIqEeq
luvp+3Qtgv3f/DGGp0ZPEzErhpz75S80LrVuswnX+Ccpc1uIfy9l5kQ0k7LuHmrceL4m3wpFO9mN
VkYqz5lnz8g1mXR8K0xoE2EYl83eEc9/N0yu3Y5DgsIxTL4fIXjx1Em6cqy1/64wkJO3WMphhC9g
SSucECaWqLtuSE5Xee+SjCzlcJXPpmqDnkpb4nAqx54aivHOMXhjXBlGdCt+qI9pkRRfQyUzGAEr
58pXZDBE0Y9mgp2P6TeQ16R2VEMDd67BPq6mhWnzIt51JvUGU+tqjKtHqzurjvxW17i8mSMMfy4H
UGfz5Y7fl4kfh9YTBrReblJd9YIexgZHTXHd4AL9na373TjDG2xRvwQ60Zc5OvTXCtHyDFNIwVOR
Nla/LjbW5l5kq0DaXtgb5Fb/EdHoLYOXfH3uFttc8ujmRct/iTO+QKasC+MdPMH1OM8CxVbccCfg
E7I1dOtKvM8vyUHZCVBzgpQlEMguz1yIKU0UJ1eYyy7fs36GjtuACs2nk1IO8/B23yD6L+EizGFk
3NVOuVU3nd3Jo3UZfEro0LPHytXZDVh9MwwhDA7+clLK9HUaNHryMRQ5vTtzUKc3WLfIgidMtjx/
O6L8Vtynggx0lkqmNa2ccmTMNuHIzYum0GkZXeN5NSV+/RhGdL0WqUMggChST2XnWRhTDTQnXJcc
jzL3RHnUeDSzi9NY8tQSXaMAQYKJucuMN/qgU4mzCOT4Ht56zP9ADbHZuII2IdOEH3pnZ0NbdXTr
AnFKNPQ7wpi+uZg9R1fjoaJkW+DVhdRVhx2V5Rj8PamohII2v3Sehwq3ICXqItkIGsWSU/6Wyf92
Ke5QrCx75AWueUxg05fPd+qfrE70YdDEBImIhwgsmATnF84G55o1LayUEoOQS+jvSEdiuS6Szqjx
AGHtpM0rnb9QAzW34meoFUf7Y5VMY4fsEEbiR4PCcolzYrwptBialudeTdB3xsGhRSKuTYrCsh0C
utGJQKTwwoLYPbVb/1AYGBqlt8c8YifU3zr5SQ4jXiT3JqSlD/I8joN21HPA96n9/HxiLzEeKJVz
/dczWIUR0xRch4FHcI1+5dlK716+C61m0fsGhWwhETXBiWj3rDFXwNkhkVVLW2XX+/XPjytU4dHm
iBdK4iI94SoBbcrP1WTpfVRnOkgUqIghiXqw6ufSHSUXIj3gIo07gEzQ/esARhLRNe0jK2LfEhIu
kNEAro64HvLVA3uOmnwkMKOF3KwzKFWJnXlyjPRwV7tL3BzgdYUzdSe7QPaJDqlKvZRjmY6woH2F
pqNW8Q2SfnM6SoFR1cLd9BGtMhEblGJFjlEYe4j820xJSw7sEt8w4T1+NCg2Kv/NF5Je5RqcJ3zD
LFI0USO+CSvjRruxjjH5dFFO8IFwXENgszn0z71Uoss9lVBAKfJydDFiICJUz7hCUZWyrS8FdGef
HaeExkNET4CVi/Q2IUcrNVAtg7KIV5pW24PwrS5qduJJHqHZsOCqrVm9HvPEubSyIYSEZ6j5Ja48
gPhK4mDSXg0lSfh9t8y0FzNjza/aB6eFq7IZaQ/57l6AGCWAs47oHw88O21thjt2/d8UQJBpHstP
wqgq6B27sWNORUdXNVB2v55UIW0yczDGDBziKizb2TtLs3Nub8Qs8AkR42qldrlPIXuDrkZ9D/0Z
C+wOmOeIcuaB14dpRmqtG7a/wmBlY6aVRkGa6XdGoYxgareMoZsvqbvmXAfJmFX1MagyPS3PuooT
lJ7kR7SD+aVNqXa0MHrDPBc40SclpN4E+w6xD1fEpkB/qe3voKSu4mBYlBkby4ytHT+IpSIJjWTW
T7xDD6j4yzap0nt1uUBZhei9Bj7wwmlu75izUcHbUPcVA07KW0VHKGFNFNcif0VBZH0odzsNWn4D
U8RDDJwo2zV8Fi52O1STyC9LkGcFTq89+Sl42JduiOInegxhNA7fH1sAcwwNPDynEqCBCnrj7pB9
mFfLqfxxEFRR4UCB0EnZDuJyEDZTYItbeUvWkLelu2hL3clTrQbOyZjE1lChcmxY5FyGxjn1wMm0
lfCbi+Ooi2CRg2glxLDTSJQ4U7FVhST4TefQHiW32O5DFsSbwDIkq7dXUAPr7EW3u1/6X60gYVMT
vcXyn2wmW5kNuTZJbqbnk7TUudzHxDR87yK7Ehdj2BDN7QL841AXqSoUc+IMLHLU7qb3rdxe+6rH
NIwjcM7OlgHLNMsaWNdinYo067i+/w8HxXx16vdUiKFA0Wnu+NaMy2NO2SvcBZHGQNtxFeB6vSBo
wsMDY/gvrnf2tuDTNJzKy7+l7avyLXLv95GZrewzu9FhXx1J+Betwdw1d72xYY6z4fOtXP6OwbfE
Eke+1JdPnZrMZqym2NQa0xyUe7aKfSxCuU7TMUA5dDES8zt1fJl58X1b6/2P6in41XGf7BB+sfBT
uhMFGLsRzN4k55rhI/SM5ckcS4wMbIPsw8dLd6wrKAHbYo0866zkUxcUqFQzHJC5aPRlgxNO3rGP
nDMUcznqDBmbI5XhCrliJ4EXz5DewbmEgV95nSb3DT8zTMu+sKaGNGPBpRUv0MFbVzn/6CPmFTeX
MFIlg3sNScdnN9Wx6Ox9W7ieP8EQIZxP9Wg6Fp3OawnBDyJ8zIfXuYDAg0idtCYtgyxxDgFBixrG
GAUkAEBQkJ4NvB6B8omaw9C+QJzbVyCl/7OSmJj0Q3Wgwd9T9LC87YMRSLml85BwJiVi3Js1Jfy/
m/UYOn6gAi5UPRjr+wXXFpYlwrv3nHBeph2yGAeBjFoLpiX70TTFcjUpS13dwq4j2vTcEocHfzPL
d21f9s2iv5peXMzb74ibnqewQDAd6epr/QpUzB6qAKdSnkb+X3bh987hZrpyjIV7yPOuQuFrhZz+
eazN0XQ/RhUVxAnejiaxwJDYe3B9hZpnp77SSfHSRKKcv6JaLNBFDfb0rhYexX9lk93y9+0sLUXE
tDndVW3Ch3Lua/K1k7bWFRy67ZP2muBlHyq38BmHoM2KoYWEjhyHEUXZtv2prEjA4fhgOePVUa5Q
UY5Q26byprtoL9A6/+PB/Htl7wyXR9nomDJPXjOxQMISfVFkFdDyZtWEBo67IuDfzzmvN+bbKIDD
Qox2CIg9Z3fc6KFfE/FtUduAfqPvUW9jNy8deWAfjJxbafzMLYefdt3VniEGyF7FVuq2eQe6jnd/
SUhHH3Q+4Ei/fc9VFAd5py2bYrxfQaPvAP7ue0vneJzshxfb7sJSaiQYcz61Y1OJrAJt5gOO2NIM
BsR6IGMB7iIcgRJQYklB7NMmDSSFYVRO/pFuxp8joxk7jG29z2lZfuqSzIhhr5NANzAReVGPa44+
pIqVP5TpavP0YWbK5t5EKHVVU44GIzG6gdbLG0W5iF8ppwx+SSqq7Qn6Lxxg1Rj0I1j6t/Fh5o1u
Ft8R5/yWpYvJgBlDufUrmVKLNq1XXyEdmdPQkt6/G8zOwZD+E9j5ShKGFheXGqXXiGwgQDlMEJWP
SAUaLQ49rJpObL/Qy84If094gjhHGjh+Und8eBmxsG2kNgLC1lptG+fWLFvQdtHLPYvLweAsFEwo
kdM60948MkRBegypLvd6yRrN7wIAd543K39Fr3129gRr1beVIqLQgEx0qCTekp5qXDkunG4S9eHN
cdPPr8kRIb4QF6dm7LisfCkOcVMS/HKl16FAf0xpK4ekfLec5TU4Q8UAh/Hy2It7bEzaMLG7ZVc0
EQFbSE8KcNGtxpR3vNZu9D8zEF0k+sU0npCx8FKdq9WDC+GU44bBMsd9tjc7yLNuJakEmGRSVMqV
GXnsRST5f13WAuLMv/iGDeSQwTwgr+q1VGgTnMmMvJENbJ6Ruo18qmHGXPgFqVnJvqHtlQzF4vH5
TT3iU85waTvaQHY0Zq1deOtBhI9NLZfLo8iGLPGPpktdIGiBvrjadomuFJ3iIQsqIJ3WjqQPwj0P
OYA9TgHNWaPZ6qKka5c8bwuMUwfQjJOppjb0zkuXE09JkWyJE8U1vgqXpkUBn2xuQPjfEpob2VmC
HqUJr5mlP9bXGkSw2aOrpOi9NXMfMUUw9oM5EJRTSZk8iI8ZVwI9sg3s6j2jEoqnmKofw0t5/jBE
1oPknHZvy4a29SpX195/37UuWrnqxR1TIqHUwLky9y2jQoBtxlGTgoL8i26FD70dD/TNsSpddDis
XZTTEzNsY/ixbFsCpCQEg+N9BTep41YHPJbQ4yQUQdzjUAfR8HNWeQQybCVNtbJqeZ/Zh+tpKh6f
ROjpNtrWx1OvQF0wG+ihtI1Ax671kao/mwZ4IaQG2U9qkxP9lvn+AYWUv6Kri1O4XUlZy7083GiX
XZqjX1XZw26pFPGkucP5uRs5N05Ya/l7pcVgCiGDJWPpcXb/ymuUPcT7HZIGPzufXOfyBj5H0whh
3qhCUFUbRa5+K4rgNpMH1u2c2kP9zUOHDH72ibqeENw6xouzoTe433kXOwjktas9VeHqn3WnKT8f
3LUPN5Q1Nq/jLsrxHGOxQYd4vlQ8V7XoYu1Phyuh6kE76R97Nbywu4/lb3kVJFkYzFgHYqi2vtbO
0tJjtWHvanAM4SxWxH2Hqc1isbH443dZbClyUWgUAup5BQh/u13hmr2tBON1MXZliHOPreljwtYP
SIpaVbkKsxPzemFrAKqrt6W+AhUSj5mR1lK6AKyQZJpAbnWW9eOonP1tiFIuaPdsTlnj/HDOvb/9
CidPNZxbV4LEnBEgqhsgBG7atooNQV1rYzcQcO2caJeG5Sm7eFeitTWm8CYTP3oh0eaOIQv7Ywzk
qeiSxaSPGkPt37+Y27rH4PFMdkLb7Sg24tC1lRqes2kCZfPEMNOhXPz1srHVe7AwcmCq5158wIq9
E8uWEo6ZHuIq/eHABfua7+h27EizkwmXlt2S0xsgFExKOSZ2BjbeoTrR4MnGyEvm2UJKd9fimELx
AAuvIWWbSjyzQET/n9sC4rlJRLh/MmWz2IyLXJNQ+Z58hmfaAbtiZfwdJplLYFP6f6eiiZuFCv+X
jidhG7I4KyO+duuDS7P8GnYAfp9Xv9RkJv+rfjmTKWF1Sd0dtf64/TdWMC4N05j1QLrx3tjbdcFP
9X8fapUzb9y3EUwTL/BXzVHdi7d6skkbB1cz/2R6SalohRd1IMha2vqxiimNFyrNON1vrFNjZWH8
Dld73RcDEpR9Xiv7JKucr5mzmxJLrMINBNwB5+/X/Oib3o9AxjfB7gi0J+TNgpxAShPPUy8vgIWw
gdZfaR6h8J6yCX2fmwWzSIT3SiAyFIQHSmzLxu4kmzfx/5zU71LWQ/kWOoSf1Sx0ZbrIVYrfNEWW
AF3L+YT2QMeT3h1kUDjvnPE2PFLqGmLLPvfB3TfKeClyG51ikMcbCGg7f9j77zbmLDyIuOqNi0Zz
8iZybNGnEIV3r50HUAgVibxOBaoMUtiqmrDhCDomph2ZmtJN9sc/EuhjuEZVy9qBG3I5MIGJe4rh
Joc6EAT1hpLVM3DbI7H+5Afyy45i5zi1ReW+v3klJFMvufAOw1JwyJU2rYRLDc4fUtafV+7w8CEL
KQPnhKlUyv7SKVHCKtDmR4qPiF5Z/NfaJZqNGzQDiGn8Qo3bIuQ96fEE/ZzWegBxbUAFJFwEnuAS
9Uy4wTqsU1FV4MZg8tM9ZO+8Nsh6LaFsEzCgcRSL5hHKG6qr28o/EQL9Ym/20zr0+rMRg6wI6GoG
WkMeHS0PVv8qfuYgcUOSe6Lz4j5+taIIF+EUcwEQwCXytjI9dkj7GZgHhyK8wWVcIvq/FmXreKBM
2aXHrnLC8fnyPnVm/yqXWtmvW4dYcBARpSjkb0pVRv/fR4weevSwpbfo68eaj7u7V3Nl0+AC7949
KI1WWrzfzMLRBrJZhslf7xx40uGpzyIrhhlnc6xcPN6ckgn7a9ArFgwoV6GhMA0bQTHkCHHigIJ3
Kg72jxvAFX78so8qe9LW2AQF9vXETALN8+zytRMuZyow1n+UEiRZALJe4a8AW/poCznYAQ9Bz3KW
GmT/MioAwDnryz6+5nelV+OvHmq6Q9z176ltqIaKn9nrNv9FnwpnEqh+uwkrSttg/oJiultN/+Va
kTPVNNQZG2cJyCLA73sduux8oHBg0s+/kJYnlBNAYuypff49FX3y/mDnok79EZDpgd59nYwy4cc/
oMtK5mTDShGXPH7wOYMBk3QvfcNhkOacvZD+x+lK0pbPQA+Sjl+/N7GARpilgjU6O10IMiQH5Upl
tgTig2XQoXEiSoEy/BUMretavZoxLeDJqt1ER4Cj3cceedGOHvzOCEq8TFShd0bnJMRi0lExTcLQ
JM6SRIjQqKbts+PuLye9NWtexylF6y5xVBsXmM66X1ncD6KVKxx8capBdwEYqKo9VFDYM5f2/zgE
JBfSU4JNUuI1WcnZW7zJ4iIRMMmSWSNi1kSmVE1PgYorSPvocvgFRN2y/SftAcedIyo3DhlK0sdh
jaS9scJmF73SfSwc2ST3NjOKmQ29+A29G97DjMzDdyx6r5SMI8eSj2E06sqroO/1Ygg8gx4tDXYo
PqSqAadftWCp1RP+GexDO+E+pGlzCpc7INW2MKPXU1hwWUaXW16TI6fKlgr0qS5Jq56MzqU5cliH
SLPTZ2S+XkWuZTxweGZSKU8HNedRLSCjX9q7WRZLWIs+lu/KF5dDDNBtPexAo9Jhct04ly8aedyU
NzVLC+k5iyiwk2XxUKnjik83JAbPDbp7wVlRAcK/7tgLy/b7bmh0YSxHL3KrwjxZwQsPV2FJLk0x
e+CDWQUDsTbmMe/QkdwiZjf6stj9hacPLxCvphJMqa4F9x57PKTc2tDFl/H+HkX7BHEIEh10qplq
Ou5MNWiydkPO/Su7IfIjKHNqDE676jZHOKRvonskDH7rY7MaFuJi1+Z/yalgBpxLoaieSBmDFG4r
HmJj8FFMp/v7lH1pn8Kzy1AsBQ8tLjtppw02ZXfCbIgjm6Wf8aWCgSlD/mSbHOagFz5UpdOXT7C3
z2+Qtn9SOUPq4ZuTHpRLCILdAEduN7cuuHed5bMGxTfNc6AmURYsvE6IDgEu8rRp6l99g2z4y4rA
D3nTe5L5fw4aKM+LBxleizv2oP1LN73DbEmH2V2c4vLBaLwDCox4rAghd3+0vvIbrxxECxwxo7Na
Vz1AylhbVP40CVxjcpmHe7d3qEAWecZkGPlFwBZh75teLgKwXuBY1FppUUu1zacdCJuztH3EoZw6
RwFnLZG2SuUofJ7zcpVHqBnggM7dE0jyl6S0owvJ4Y7/I9ttJSIIGXjaVJ/nGPcp71yR4FBt2+Gs
1mo4qsg1cE+41f/lcR/XlZANtgJWNCRLGbKTOLRI3CZtLAQQHN1aQ+wPbieG4ACXA4+Y+xJ1y7zH
PqucMxFt9bsWOB0VaG6WQgatPKdn8dqnWgw9F1sPXi/vDqH6reIBoIEWVOg0XE47cH1y5GZri6E3
42pnpNQXESWtfm4mEAwBlwfhepAWcrIFJXYOtwE1WDMvUom1JirF2d8NYkaGvc3m+WXu6Y1xRNur
l+g0VkKoC3nCbBeLn7J/h6Xk98U4QLLr44IUuteNTBqBBSYDnD8jlQm9MQcYypSZ5XzZNtQd/Eyv
E5+vnsOfJ0FV9TDwOgTZxv+pWPwGaiRKpkdHr2yqzwtwHSSA1cyvG81DRIC8rwr7QV9J5+YbDm1J
zfA5bWZNhqw8Dajr0qxXEL+oZOWMQ93tN8qFKQHloGz21u30ScUi10awBYTeh7q5d5SnZ9tuRprW
y2wprsl6SXjcyBLTLlVir0bhke7YS2P98WYzLgVBjt2MNzrNJa9XB+OfrGH+CmJ8ypeS24NRCyFM
l0GPNZ/4JUZvgKx6FkLT5AujC7DA+tKV22iEOrAWygFAMSZGA70C9Cx06j7ETYLvB+0tbPVstJ+C
d6htXbq1DEKF537gtxXwhvYGTgPrHce+GHyLiQ5xHimo/tU9j42tTQg5pUb1EaeT6YCvoJYfk7hl
ow7Zq5avtpJvSKH9pfX0Uv3i+qlF420fVR2wQ42BZ2F/JkfJoXRsQNz/RSErFVO3PxFAU+pRkxgr
d6oGXoLNtskFm70YeZKh7ezv0nywv3jKbY33ShxRhqixxLnIF+nmM24kflYLzO5Oj28N7Xl7N8AF
QYyWksfjk8VlXwrUle4XeDfFn2QK/Uw+B+Bfctg5QRDzLm/13ylrUg6cCb/4VcxTg7dYbeUEZIyl
nFlThVp5XA3hqWJrz1EGnmQGcvzjL6TplMQlCka4VhNqHoQT0rW/99egq1/iGarM5C0kNb2fZoQG
9HxJXBn0urXFDyUCKPbYzi/YJpGV+C3zG8Sr1muw5duaMLklv9lLczguMr85fBx7P0TSf4KDtSYH
VROu6oZmnVU6lHTcYCgPG+jqRLxSD+3Jgmxud4V9gaaeunrYLg5CVm7rYlo+m5Y9htkdMFAu0B5s
M6QR6/stwHn7dA+N5DDHN1tLnBfIPO4tLPqtHejQSaawRYcGx97Ed13sClMLBaP2FWdyGDmoCZVO
yeTHE8aX5JLDMYH/uwsc/ltXsnCPzu0RGFEaiCtbl0YI+NRYKVVPPmkDiA6DniTzrF80i4q/iFtE
ywvyJDirNuBI/Jfwe/QRaIZhfbeiEFieXi+JjsLNZu+Yd98hMwxd4he8JPKZCDWG4TUPjw4bc5U/
pf5IjN8Qe+tQQIExD9ZBdpphXntz9VY3CnBWPvvFSqYlKbDWnnuJnnbjl2h0+q7TDtAxYv4WpntV
p973rLfWr50auhk8MKPRIDW1/nG8ZDLksZkVmlzhf+iT6wPIhmk3xpw94rqmmqJBOrqFmnCltY39
JKHhOMQdltC/IR3J+CxxKcBot+9I/qjKvcPtoxSOGAQcELDBxS4hPdre2x2LWCk0L2uR6CwAiuuG
S2UZSRZxLnk7z+5XubAqWxD4v5dSQrBW/avp5UFPLAqt7zzCyx5LkmpkWwqAuvoNY6SMCQYyDyH+
t8sKlSViyH9C1UNAketwZdQV/EQNz8FUrgSvt1HlfDXSFfC9SGTQOeGLfVtyPMSJSxKRj8rjY0jb
LYvmoDHEcUacDi3hDOMgv9ePVGF1tL18HYsLfTsh5hGgJW4v/ZU2PIfShxVTbh/2ux3joaiJFkaM
BciSRUWmXsvdY0EYZ2jkKx/LAvyIlnp3KtHyKeXVAU+cSyt9eDgG8k1VU1haOMBmuEAVUkjIH037
ukngWxIHvfUbSNNJfW5mwkpJ73SaU2RJ/x2XKBIOqBxKQx9PGwBb3UhuMcgFC4T3Bgef2tlK1CNZ
6rmQe5eCBt8ujS0sJiJdehCVrhxDS9syCVJZqLvKx/fpFSxdNOABsOs2xb+TuCp0SPsl30bQrKeV
X6o9RfQYpLq1gicthJPbiCH6/ArDcsKmoGb0aSr2I5G2arzLw9cYpkb9iNhi3tS6PcuDvfqAerIX
JMA8uABQVF/UwfzAWdUGzgYpEsLUfMRPS/e5a4nhs4YcJ80A9mwGucEYC9LNxrAHhr0Y3C3a8r9j
wx7yQFXwGtzXVOCBi4zHhtxzCnw4M7OGXVVgAkH+PkR1JxdBo47mHXP83l7ZY8y+fIBxVmTBN1kY
Qm+bCVGf+Bdgi8AxlqTCvZcFPuZqhQme/prnQ8fhg4BiYT4sgns5EeVfStIDHM2o9I3IKh/6n4eJ
HtML5+CV9p9+oSQJrpj7Oga3ABOjl/UfxC9TCe3SO0HZn1BkpNG9/LhFPS8ZZ2Ia2vsZRtN++g4l
HzfJBaW6Js6aW4d+/gOTUK4skRKuLZnC0xO6iL/ReB+CIbeUUHNd4KlEfuX8edLap/znR1QcY2qk
7ftcef0y3ayCfDpZfbhO91W3WTEgTl/+8Nlag8MyW+kQ90VKN9CmjA5TngnZOZ1ZZZ9fe1N74Q1/
qHpEqFxuHFhcDsj42WHHFovnanqE8wCuLcPHapDFyaJPzh+pdNLoKIR1D8oit7w9DYt7H5NMZtRT
RGCe/AzhnbrYpTPkDsybS865UsmsCN52fHom1lzun7vcpmUK5N8Bl8t915sPVUGehe5Rce/WuWmJ
lMUcSKqB1obrprOnxKsBsy9TfaTZIIYdOpOv/KdIFMFSEyMa+aUODTtha49H9S5jNs958xS3EXx3
6Mmdgjqr4L9wYubeJwh+NPgsnDGJbmvTHdUS23DADao7ZhF5tFJ4SIm75XFohp7l0x9DFcrQUUOK
AL5Z73Emy6a95CPOfwq3Py6yble5GqYM6h4DXHFTPcY0Rh2z3RsTrTEVrai44AgxuXQuxiJ2P4VJ
b3FHjeiKZgL8czxpFA9B9wBgrAycwlljhADPtDb7s9Smx89SPx396qTSMjIa8WTMY9A0Clq/7bfd
/YrLdAFPrWtmuB+UXZeQe3JAiMoZaUiIZpUAkw/FMoWr49KklKxY1Ggz8xWoo9uQGnYzLiOktwl9
g7Kb7IMxgMHqhxajoEsPAeiDk/sDt2c2WPlmzv28QDDIXH2QlGhn6HNUNGj3zf8r8DLa2MK9Fn75
eR6I8RfVeBt+lyv4zWYjxfNiNQYcLha9+TKGXNbf2wPHavAYynyzsbKxmHHdJayacBY3/W89V+uQ
zyDnVaIRgko5InE5k8M68Tl1m12Yon6xVjUvYzXh0DvpZ0aTL0Vg2p+kzsYazKyA8ejc+M9pFZDD
/MeayF4LuQ89VhqdlOYTKHqHp9IM4kJumiLMhFaoIcDk2kVR1131ps1Dfkvr8Djqso4oZbd+9sz9
eDOxz5crhc+2bJuqeVgjksmK2fJVCnOgaMNALWyrifA0wm4pdsj/Q4K0T2PuvXvAy/s/Rqo4gYOc
466SnYD0FEyaN8CxO43WKtDNakiho8EcY/Qg+ohAgkulz2SwUxOok5vza6YHXtnCvGz4O6rZEXv4
seb4RxC8WQjvDOiIQsflGIt7ZNA+VhqTqVLCuF08ReZ+3xKBI5SS2ZutBRcSSQSIjyRdMr+RRtGW
l71xw6tHVXnEfpntlPv4q1CUxJa3M33DRiUfZmtbRi8obckn9uOa6Piqo90QTMAr7o9VUqZb2Wc2
lwlEbrwlaYG+BYq47pcBSS5d0152SR7m5NpieIG2K1vABnTvrwR+WQVL93z+H2iIceZlwQgGOXrd
lF5b0j5F2ijJMIUarejdZU4sBjvWXK89Bd/Nxcor2xlHEsousgI4ny+/hKvSENaL0It5ZYWnL3v1
ZNU/YBKg544l/pcjlcJ6L3dvRgFQWy6oICLwkmi+PsYfuJUZxxxQWCZWnKq9JbPvUkD4KiHcdcrO
Fv+W47FgjJ/DIgyK8dxO+a1VLwR6//i8PtfpNI8IPpCerCENOuTrNAxy4xugG3MPZbqGDJT0lakZ
02aJ/ICNVRi+/FW7wrKdkJ/TGjeuatvviDTMKiRAygHP87KcuWQ0Az5tLFS3WLs9sWxdNmgelDi7
AQkthCrkQg7SHVvXD+UB/4ZYSvyPbk0fTmX5ZZedivFADTgxVOAaTbhrrt+Bn9m+cEt67A/Y88aC
A6jN9LogzmFQ3oFaZhL2zNTU7k/TGC6v8v238rYJE5640pv4ym5Fx++fjOHVmnZdFEzG0xzw0O3S
41EiJMIft01cbeCDXWk3kk6gr7ogB0IdYJkghVLJeUmrozGrwnQ1kyp+NAORA9T0Tb7JF7WEjLL0
awQpdkRt1N9CX6LVxJPZE9jB09auUHIS3k7Cdxmnmk40qe2uMA87udxFUqiKi4Ox+xRz8NfeDtIt
rkX9st2EW9yMxrqDcPcL8klb7GjOroFVqy+Lt5GNI2yIli5tp5A0pFY4AVHSd6NJX6D71q+/2h5C
s6J1JG9+VO6Jr7AK4Q6KoXtD8/0+WXwAwPKT7dFZwnJX06V2TtS2SQNAV+xH9eIvcj1a3QW+BxPK
JmpD8f+FDVnTYHxNQy0Xehl3BJabac5pdYNDCBgMumrBsKU5FzdKJErMRMpz2qRBAHjvsFl2Wve+
rtV9yvg4b2sn2DSeVuXQbR1+ezCOKQcbrRFltEriO9T0ZkTvCuTGZt0daJv57ahW7SLbomhz40aV
/jxmtDEtilVgIPnF6jmcXxODJSQ2IxLag0vNQdgYJmW4Vy6yoSEsI70EVArjIYCII8sGdy1pANJG
nM93ZtyzyV95DvLfvuiYhaEhHkWF2ofcQnrAPY5HLl+i/7djIUFh5oVQlLjAduiQSKIytgAUCDDZ
f9eBK/l/C89VfM5KAeVf7HpiD+ZC85l2yOgBZvv4inO9AEsYWNev9N1J25Eu+h0jUYDt52pmya8S
roUVVSPGLVThdDvGgtyd54bMZt9gGGNWM9U6VtzatzwWwJmvHuZtkIoLuVbJDe7aNcBn4ZM8xUpM
S8anmRRLVENgfQ+H8/uVKFtY0V4wmk6lpe6wGFE8fPe0vR8BxdrTCuIxa3e2Yh/T4BIuKRV0OBPz
1LFbJvQ21x7tq9b9gNbu/LTXb+ZKZgbzCDLVbl93m6x3aUWQebQesN8zeVG5xpLrV6o/86v0g+Vi
8m+DnrkFLZotA5KbkjXCcsZ8qZaUIo68KauXoPOebK7V/6T6bxE4vP0/LkYQyVuwWcc2IHdixF50
xQM5YmeJRbS+haSv32PX7gUMuhrIytW7RflbgfXxahTpVCue5+5vqfIe4Aj6cgDov9KrKkhuLLvY
7jjjzZ3oiYkWa1pjGjTwrrWiHeK3dr7cl1WvQ3e/LX1zTshxOfBvu54cw4h7GaD8JnJ8AsQWnu27
wEWA9qg8HpoKZg8SfzUwFLVj7pBrav9ljiTRRiwKeticVueBAgG4V8z8/xgcsHVeZN+WJEMGSnZI
0HczrqDw85Yf8sqQ6RweFnjJo2cU8oBgCTx0oz/Pdz11gndoB1bZr9s7ahT2tXWeDkLXfNWfoqvb
Uc7rZVqdFwy/yHLNgN6bW3uSRKqBVPdAOL1ljEizvafylJQtelWqbgQZzY2p0j8wkrRoW7Bhfnuw
16klH/Ha+bp0qcyNcdp/OEOqf/nnbW0/x8wjy4PBGR2xaHhlhGoh0BFdrm7nxDNoaO1+I2kv2ibS
GwSOEhqnE0w4t25yO9XZ5alPY1sowStQG8f7AmOYyHYAdQQPR1pDAaxFBqmZBBxNYhOzntnKevfA
/rhJVH4SpHdvrWpgPtaLg0Lvw3VkSsSpMthpEM4aL9Qkdyq4C0D6FfwKY5mZUUzu5f8BCLvWQibt
CJPQUYz4sssaTql1vAeTaNzDwsnhv6hZidTfeud7s7BG4UEdHnuv5p3FDvCzeDSNfykLo5iYYSoQ
/UgtBtPUBjTh0Ua6rWmE/xXW/jeErFj9oYPyTDxAU77Tvuv7P7vkNRiEa73hDtTvuuodt8cKfbfS
RPWeFDcRn+xg7Rlrdgke4aoVAPvACZQElyQ5kFfmtINaqf8IIDbjxEOL6O0xi+vyRj0f39n2BfJs
h9Vx61QQaXvqqsKRFZPl73d2eHLFnGOvZBLTd1vGfZD1LuEupnrIhsbBMuEMflhO5uiY2+/6Hd0n
dccjnN4gFOqgZ8PW4KyWN1Xjmcs6rt5r1GncxFiKuu/6TvXihan7XuMyeis4abF22epdSv7SCZZ3
xyZ/qx8PXXj4YN4rpwrobJHERgLydambsOtZWA6ANDUwjjNCRNHK+bF9L3aWs+2YJbPecdhuNr9B
a46Yiz4T8S+DHj+hswzajLZn0ME5hfaVD+Ec0E4h/2LgeWzUGSaiEyHdhg5cd+ESJ7NzcFwaOWlC
1kBYQzSYBvbFpfSRhzLEV9muUf7mGmIPgxzZER2gUq3BF9Ub91BYYTee9fs2hxoVyapqmY3cqEVo
ImW0ngoDo2qeJza1xFj2Dzx/amghmEK5DPweQhHTcLCiEXXzDnyL540HkIz22lO0wD94HwuhP1j6
3dj+6a948Qt6zEQ79xPUAUcBlLKl2robHCuktunsY7sHAAMiXRJGTHTMj1Ka5U+VTS3tKWY+2ujF
QlWLT+DO2YJyAPi9XQzqu6sEQmw5CRGjcikOsEjjXXH20mKGI3WSDbJ9IOeKGMYjEoRktyQrTC4b
FmTut/4wHcPovZmPGkxlX4zg+CWB7dnsxEkYy4yunQc0FvxHQWEne8fklYcV45iMSBKWN/H6vLTR
kqTFo9GdfiVV8J0KZLbvF+eFhCw4Btp7sSX/0sZk5F6/7jbro2q0JN+KDDuKoBXt6xlUGNKl80Y6
bnJVSBmewtoITji18snlja1XVOtmcBVQD0zTW3DWzzof7h8+RYO9wCzev8b+beYEGkd8LrKar5O9
uU0dYx4oZjOsxGV9sBBQEGGNo60+LAQCSa00N+whf1dPEtrNgH3noF7du9CTGMpwRGjIcOhhEV1I
kXPVulKlQVU+wJEXV8szaiuVbYCSKZCvTiSkTy/wsTx/HbMPhrNWmzTrNVTfDiymn9PstYAmhmYf
ycKdlKtMdpJhZ4IU/WA3Bji8Xc4wU6V5GtqjGa/uMFfrfL4XfGexqf0Tr1s1BuFEErTHot4TTTZ6
A9kGOd3VSRLbO7re1cV3E94FvlUlA7n2DoZbns3YXvyA9wbDtX1uJv2mmQMVHCUwWNiFoLucK2DT
Ha0UgKaczxMMhpReEv4fkrAqBNonybBbABvgA+SdhQ0xYyhZHQSTIcBI7KfsevMlWDIb7QFhAOwT
4xmp2U4NsMNbpz7OKSAbG0O76gKQQE569KY5k54aIEN1luObMMM3lcyyqjJ71B5qW1gD9Zn/rCgQ
fwsAVPCuddWkMrPsGFylHGS1GbJJ/vqqM6ArQZjKt4C5q2eIhK5DLmvNUee+UBZ/RgE8YTUfif/P
hR7F3WiOSioE3fEDWRuCJvbLRGnaeXwpGgXpqDeG2T4jW3mwYeOBtn1auMHcPupcH8OyFdiw7vIB
TaHa8kFUCw3sHvW7cWPDzFUvd6Fx4R2WtJz/sArRIYucJhLvzVsi7YDbCGZvmt4lV2LOemkw6hP8
2EeXCjgNZqIgfGS+gUad6jcpWhUt3HQNpxpUCz5LhMWCP5MQbQlkaIq2jIksaoJ8vp9qIJ4DqxU6
+HkLFYiPxBIwyrhwV6Pr57v6nvDR9jfS/Z/LGWBE77QhinKAbSY0AHNyMVGZRm5+N0R3TvZoAL+t
P9FfZmmY7CW639CzoTErHTwJWVtja32WP3z3aa9/zy4RtzYVblNBRyeZd+dsjBi7jsXh047coe4h
L1sDTXWKFSWCsNZDIZoSmZiFjUSukmHBM2dnYJrjWbl15UxWZfWtXMWop0jxCYdPKanEbU8DGiAG
1OGPUOoOv4Rkefa9iwtwkgcqvlopnt/Edbau71Q4fYljGzuYrJIhDmew5YbNi2/DIpikyB9SWtWB
qujQtoAWFqJpSkpbeh1P8hthgRhJP7yMGogN9etJtoZObgiwlErg38ewCWwHqa5nc6lbwSUseZ+e
JZdf2Jd/oZwCHFzO8rex2AMdzyoG9sySZUmhSP4ZTdipnR8zaQBcocBvXizR5Aau8CxvBKXs7/2J
/GL0qLAZkagFp/xBBIUFwbgXou3sfpiE6JwCyaU24cgtzcpbJAtDZVo0ewhS1z+6YLzL0MI29i8O
GALSkAHBB1nZCzx/0fsAdwFXYsHWe1VxdpP+SKNWYl/uqEdI3MjAVx00rDeAc9lfcDsvIwYuv2Lu
x9IoUqHeUxbqg7Z26AqxntdYbTuMFCrJcLDkK7ttZEhy+A8oVOrg2yIc0iYpPG1MNAzdi1g1a6SX
SJDdNaByfjSQcvsUWqmu4nUk54sG66Y0vPdB4Cjhxf/rQZFP+h5PT/fKsAgY4QL5342TL0IwEyxE
pL1LoG/zzRAMif45jg17HbT0WWEsUh7y9AxAkgJ9LFtIgLFfOML37Gc8HGxfIkXlOB/d9fnAA2cH
wU7ZrBJCWKfCLjWU1Bx3NEwF5If98l3hRWS8ldTl8cBZlYb4jeGUiCSerOUR6uqAz+C3TrCRjqu4
sgMxTXpBQOiFn8FMLSjirbOpPo3MeQISFPkeMPnYIcip9q9SORKhtkBinDCFF4NxhS0adtW7GZbo
bF+88JZvif8IqGqLeEnPxBmQ0AKGwjqvyB44S0Mbe2ulr10d4ArOCvPpFEus7/nKQXm4paUB64og
+/XoxJM8u0xGM04CE8rEwAyGzZQMjHQqqkPPMtnIKxZTZFkKUC+yJMnyUmx2bU2LFO2KunlP4JCa
k9ipyrPChOERWxaMWHDauBOmVy6wevXEv4alNGIMvZbFGn2lYfzIdToFDORdITWsz06f0+LufpMx
4pkZdhbxg+NShb4FCXyLru+fT1NvwReiOZ0OhE2uaEjSDQ1lNR5uSwi2L0boHliXtQ5mdbSjjKlS
UE+2PxbTzEvIlq3s9uwOlQYA4HPI/Chh8esk/3gvm+alFdgN+ZkjYG64jkPpja9ZQUDygwFAN4ia
4Ukh42OAfk6wuVOof8TawmLBYrSpOhuU/dR2P7rwG9EkeBWbaF7zzLXMLF8kcwSNE4BE5IgtUKlP
uHPhF40h1pduwgP4CuUYUbuEs9nIRAMs9Wp8Jeu7lZ5yygZ/CtqsReDwrdNStI7ZQwo61LLAIKQq
3TZEkyG7xIqzUhW7P+zsNlTLSq2tJ++gWZw0mTQ1IsXHW/YrSDJtAoDnDj3WO5UksmLZGDXtQZ/o
Zr9+p4k6AYRB3mQhDLGUCAKa0etdITRHNrNoNBOaeVTAhz8YpkwPEo4Hb5XQUlpR+NrkxUBQUDx0
4ylVvDnDbF4Rmx9n/ZBNpBeXm+VRBVxbYhJk2Ggbs39ydk5DBUu3TcS7tVVUWrzcOA/91XnedqV0
KRmuXMR2r2W8KWt136vhXsbAeDC9LiRJ8sQJcTmluy2wzwre+FdLJicIKezyM4in0u5MYXvGMdDk
xKsempJwfzJ4lZP8wAcrmDR8wM1WEvkNHucGuev5+L9lQw+yYhZ4PreQHr5oPTsNABsUFsc9Z6eS
Iz+828fja9MP0+Jazqofxx1kiWsMpttIdeMCx5/amiZobfPdrlEJlrykXgNt+XheC09iAQ07H9R4
dzBVSv/8ycmsOTe4ho+GVtqcY+gZq7xM+Kzfx1lKUnfdh+SYC96UxZo0gHm1FebRFTipS8/vQqDK
pfDTF7BUuqLclqujjocJSDGTKplJGdkVOh3PUiRq4dps8+2pH8wV2LNSGTQs+qrliSvWPZwQkopw
vYG9+KIjHxPmjeBad12ar35nvdPwyOqdrfmaTgmwG672LWoztFBMcZNKUDFuOKPsQ85/RB1GtYVa
jc7nhjr7GDWGB7U20JqnFS8GRdGYkfnL0dRlHVGMaU4Avedg8tBxt4nO7dTrx94bkibbvh2lSI9A
HaUspFsnzD6P40wWb5/QZlYIqzrxfX24egUeliQbmiKmrjtKxhTRupqUgFqgNYbKed/O5rxr8Ye0
BM/Ye19u7LEEqNTmeyIYldal59aMCxQawCBmrzXomYjkIOwvoLa6fNb0dYKO+HljdRK4dptpY/dA
mucMdDdbTs70hfHI1oMKjxCbZLF2BEcEpVQRY2O3ezO7YbUtaKXSBX8w0qxQG507qabAOlkB0yJv
6aD/ddG9uDxr4ZOFBf5Ib4aYurOMXwsIhqICLRRW7q4Et9E+M6bh648xC+VG399LD96a1Z8r4T3g
3AfBIihqZzI88f6zz1lj9xdKwvWCffKjsHH3kmMtqGFgdbC/MvsPgetIT5U496P3Xy/5oBg0deTG
sXMU0Cj0cY031bEg6+7yU6CjxRKmJ6Qtw3csHgvw/C3RdSaMTgVYOJLAV4/f2/FXSV6A2O54ptcd
3wDJNVSOEdVh0fHMnDMzmZZOmIJ3Eeci6z4ysuAjhRzSY0bzfVYHZ/EUphnRN0+1Gxp56nLIZQOz
YdD6a94TyvwyvAWRGCf7QA3fpBbAErX5AZzUq5YLDTn3A4WXzeNS08fG94IiuyJZOyzjekHLl4fn
m2ZMoTl+ZmffLMRJrtG7/JIVzO324/NuKxF6QBTq7RzLmVllpGHVR1MQRth9gh7hfz0dS1NGbIda
WFiUEwN3RufIwXUxxXg88hX7NFVWQVw1uqQgGOH6M56rBs+jfcD4xEejZYozEv9+qHRvd2RbTV/W
2Di6H4sbzmw0kfdB+H5wbKEmZy0v8Y5J9Jzn0Q6iat3VE6GLtS+2uL+NDgx8jltceJFdL6A3gtcs
iM3/ALxX6UJbyJx4xAxYA3Xw52HoExFS8bBTsp2vKtfrjRiIn8EHRUQwhNxbUproP18nxnOsoW0c
ZkHn0GzAZWaq+MI9SwyQquOBhxURIh8PPaj2jvUkBeqmEYo5/VGlANl4GrjFm+ja6ZoUMpAfvjOh
Pn3DM8eO9IlnV2MlzDvv36BZkKyH9GtuESgy74HJMsd9IoPq1t8FtALBFOzsY1Zuj1fWR9gjMgn9
Kpd7QMfwON5mLU00p1SOtUBPlTG48zdMKnf6x6/+Ex6Qw4NBa6o0AKT8xI+VBg4O6ClqmFApylPC
apve2/o7esR8K8Isjh6LjUco2x5pMUzHPIYywdHPyMl/VNdBs3ZmW/UceYtQUckU9X2oExsESZmJ
n69nJMMpvXIelz+zwk/q0RFkGHJD7j/qkkjvJ/rNadWe2RVO1oFVhZG5BIBfdaxKka7XZB96EphV
6pjZAB4Q8YF4xHzQsTQmsBK3jspsD2fg94IHVSo2oO8d8KeSmqzXkf/195WvsCWdQCcKXTXby7iB
92lpZZxqH00sqmGMrQbs9omdIrWTpQ74A3Bh1vJwWPYDwSmFnJjuGXOlSHD4T0//J7u2xCWgLfeM
qMryPDpghLzfM/9hbqj8iQ/FhXg0XdRyPAL1UTm8GfMs42nMya08v+3O28CbrVPVRCW3YswDi8+l
mueK3IAlFK9MYJC23XhsJVqfp8f3N4O/rLRxTPXYxWSJs1PG3o3sJx8023UkibKFLRcpjK2UFAkY
Z0kY81gKuboOolVtUzJsrzBKiHW6ZsT/TebTX1gICHGITCAp7/pzbhSW/CpqwYRtywoBqDIo3Ej6
i+JS/3/+InmLfG3J0WNCd8o9gIUiO0292v6x3DwEHZmAGwjJ9ZILnxZz59yKz5Y4ozhb44kbPJqK
RmDPiZkxImlCQ+jH8nWQpaACUvrC2dBRwkxw1Il+nxCAEj8WHVThGWfetcxifPy1TT0ZUOM3UrhY
z3Bh10cr3y8TzH7REQPwcRtR85DeSSPbYgJg8VsSPqlTNoMALxCIZjXxV2sV6sEEx9El8Z9fZiUk
bTuZ+fEvpphztXRpjbHAuVkOVKM8scX2Ao7Cd0EeciIxfiQ3PNdXwsBUtPxDYpM7ZOo67lUDOten
qub9PNyadcKmB38Pk81fFw3j7T74vYOpqtfl7gfcW3Zv8CtkaS4aweiwih3pngawfmH06KOlU+O5
Mq7Km8Yoiq1a3ux0i7dInKyJA4XDv68CRkgqbchen+bVE/suABHO6gpwioBna8PtHeVbAQx82FH9
daOYHfthwCSkXC1RMGr/bcI9ksOV5x3vy/HVEQl3ZwlZgLhYVk/P3YpdMvcg+CCf2KLEP+/nzF3j
9Zgipt3IqHtGX5JoxrEh6nF2+g89KL/7bfDH0bpE5mVOHUBPzmQd7EWCAKu6YABb6LGjqL3ZoPvM
0Tnz9NKqeEwJLdRh8I4e12UhInX/FRs8bwCol+9XYuMwc79VVPhtyCbgqCbHo/nu2b+Yx6im9DET
kXjkFE5RkAykQ9kcEixhDZhiLXJ1HzhC5+AEAjyGsYbGqZJX4drZiFp8NU2RAWKA5SzzGhLbQlgF
vLQF06RRvILjlbdc0ZeFOcz4toE8sARoJB5FJ9mRpgH/Z+oAiWNEqcrZAKrPthdU6Wc4smCZZrKX
3wHZwWp8YeHNcnDwqPkrx3EfP5Woa8cL/AgLZ/2ria+MSZkJQZSO+YIj4pTGJqB4bSorGZIAY22U
5UgBxBbs6q2sbHSw8q3uGI6jugVf3bBm0p22xfIR+O8yC6TCXzCna4AIBFmlTelIN1355P7lwJtR
A+eR61pn8TTG7CsCuGangdy85x1qpOReCSpsjJ2C6mlLdMdWxq3HAD2gsR1gt06xbvthUS+U5o2S
Yq/ERZ3+yklWB1n42KuPis4I2QFPHIBxo1GXMEOdr4cg77xAy/26abcOjDwA50x3AcsrQIjZA5H0
lpXxqK0nZq9dihuK8mv8Flsrr93WAeBfJsxD7KKK4ozwAM1Xa40kaZgqryqWlBl7bJNg33PFCKZt
6wMrFbeQXr8UBl3YSJntUbptQJSVgdFvWexUzxffW57rg2jHV0rLiy8CtKsfcP19TGGFJuytqO9T
lhHuoAakjuu5rFrJOmF//cwnE9o+0busk/JPDaJ79SEZzqpuM1oS79fyfo/Auq/5YV/2FuRJPzYs
N35VUGx6kFnuWvg0TWIip2Rbbb8AB0wGrwFrNQp+WvhiaJjb844Qocose61rorAKD03hxNd5l7+t
G1XezjDDby8lro25rxowqejdHM2/kIsauy8lk4Mog9DIkxTTNIKOxM5IlqlhGxDVDQwMlCBXYJGj
tq986Ux7KWj0yWjf8Bed1z785IHwCHboXXCp7a26P1MwwrixWiRFJ9IU7fGwe1AoQdvcQ/GvJllR
HI2aqS7XtYnx95sVWbZsmiuVzrj5NaQISF6cGYlqIu9L3VxT7mVvW+8228rbYwX/69CLiM2j2un0
SUgQA7tyOSUqJ/1TNq+6p/Xg1hB1p7C3aRrGwyS1+qNNIndIqsXSyA+vttEXP0FMkoYRJZGxn3EX
wRQNYi1RrgJVGiH1JhP4fuEmDTCeavI//sMxC9NfrfYnQdIJ3HqiQ4jxPJUs9VibW6sxn3dMQms/
fK1L1BFrRYlnrl5AvdbNW/L+6Fn+sL12SOPMJhLHOKd+hDXrBHoNl5diXcBlffpHZhr6qnq5BjoW
4rd1IM9caRqlJRkejOK8sdddsEyej4egVTU4R+fXc5dsvmMv6H6LJHmb8Lgdmk3sUMZ/CaY5WgeH
ZoKdUQV6Z0jjpOYbqq4KKI4mPRG/tPxEJh8qe8qbD88NBzPurKXXlLuYn6F2PWSUWk5CHUq0E2yb
9P7uLVX/PJ8iUIdbNt/4pgd5RcFcIReStx6a4k2r/2TOx1YywWyJ+Bg/j77MCuXJwSat7CCjjFyA
buXCXcOsQZMsbZvnyJl+Lgq8mXQDVxm0JjqrrKUuca4L46gja4IkksdgDGDr61COQIz9WqvOXOuf
9AdlZ33jUAwJ/i9nAGwMW87ywZU/Tun4qIZxiC1brMcNukGYavCwyIOU6YmG4nd6BymP3WuzVv4A
MS2DyFN+eJRti8XAVEOvlh08iTC7QNOwbryEVR6RzniT7hLVC5BoU8YuXaMnHuroagSYyuh3ig79
We+NuaooVB6ljW0OVO7dF5XTZDYn+LeFoF407SlJw5tue5xQkwI2JhWOh5pUXqk9YpRnRwQ9NPI+
MpZvg5hE3PiUU9RwItnn1SYYito5BC8n3hrvLqbcEVjPx9yTSGW8DvKsrpw+J7ZbKn4p2vRWVjDh
7qiOvIvTLfs8LcNQj3wKslMV+Jy2YqA2emFw2o8chPKvNoE9B4SjSpqT8n8rPbzjLZJH6hx43fB0
IWJ32KOLXs5/C99SqG1GqZ1Rx82U5qhP7Dn4mA5CgnlAWD/li6xfiPCD/uZI7IJcuNwCKgWMf9Hc
S/Y8jp6zenApR5jupnvlFTqgiFDnPGd3Vv0ECFXnB6vb3A85TIX17t2fuh+zzzdaZgV7Cf1ouAKo
iZtcKtyrQvrhuVzxqYnt1lOaOoKQF1w7Kvy9EXwv8S6SSl+GmCjp7N2iAKjSxFWuu4AbexbttRpp
6xqhDv9in5k8RDsvtlHEsxaQqYNhtuEPNLS7Fzlaaq5Wzfyxq1PVTYuMgcK0Se2Z/vstEmaLEMJ8
X3VIeH7wHvuwqOwQhUeHSUphi03OKMUvLVjziTMMcpOAAQKMRwdZc8r7SP5fH98WvUdVvZlB9yRy
l9RanjqNEQGlG1oWF0+S0ef/DjCp/b/YetimhbEwsWxDbh+zKGzFX7KOlxSEw+O4A4Jcs+roFITQ
KmUzJXO5dpENhLlV81Hr4gQ00tqvTXrIueDW53Rlu5KL2Yf8739MEfmdyaJObnSaUin3QS2Jz/fr
k7xgHX+pOXFOu/W4T5LLaVjsrH5XS2sNca1xih+qNRWiQmVRGTpvkQSNNwFL+tx6382bRfo6nbYN
qyKWKWL1LyCuGmkdUdFwC59j9GWxU8d5b7JtDERBwRHmQ/NT8tBzPJ0XxWOLAAqMrEQsY9OiVHW4
KWuD0pAzjg15LqxaxTWe9YUsB/Dt/AEsnrbk+pVYXfGMK/ZlFOYneGHZZD1yv2ethnEtYVq1AHt4
26kqz6CN57yCwEb92YpGXLgw8yHHsDdCZQH7ibbVUvvTBYbQ4rApgtqLvL9SV1XCL2Ijw14caMyg
OUP76kKX+3E3K/k7onM3WUpNh6USAyM28qO/YqwJKINtpCf7YEcI6OKCvbhplh9EfBYaALUWCg6R
zPjt7kLlJTIVsJdBy8fQjdwBXg15sF6UnKDFEeHDC8MATbbYeYfLUx7kB2ZmaflJhLG7IXMw7NwN
Cg7sK5VWo/6N26yqXWyXPy1e6YF0ZMRcFtZqHcmy6++3mbQgUfvUe+g0cN0Tvao9m8XZ+Gt8HkG4
J4TX55dZOmZ8ddFVDNOWcU4lpoMZKAFGlDXRggLrTomm5bQTEkQN0A9/G62e9fTBAj5+gEu17+ys
V0w6j/kVcQsBpJHiMks9lF8LqUxL0u4ii1ZAFl8w4cHZzOOgHWDvbX2e8CmLw5ucR5QyOaufpOXn
x7t3Ah/NqIYibnTr36HCtqm2L/Z0Um6usCbsBS3NhYDFUsG0vTP+6wOTH8KkOVFZdKgQUokXTuT1
iG/A4Akz1LzeGZ0mdtcJDPCvMd0vGmGdYFaJ2eqDHNSE7uw5e+FU9jAcu1HupuY0Rv5AlbZETIH4
uIUA2nUaRTvwxddXuUK8nNmvmwf3ArkFeSRUNsKSLcNQuIy1onc8l1KdS/ZL53+ju+KBol9XcLkG
Azqr2PiaS1pSCWxjoiGLZAKDbbCNZz1XR05TJF5DO7Lm8WP+pc+81V72PRaDv8SMmfBIMfEunRzF
rSrOkp5b7u7dOuimXKjOKe5g/IQsLUvjz/YrnUIP4bGs8WtQFBmZscw6smftQcJP8pbjkzahgHek
ooak3NKoxNAOfV49e3aPH901Sy7n1KxEAtp1pTj/j5UYEyNLLAHZVcuBvgN+IONpse1YbL0sgQh8
h2DkpJk55xNq9UqjbtIYNiMskA1qvahbq9IPokzBKD1oKz47YbvuCHQQFTpfauqsCHLiJ1mKYzBS
NyNtTXApic9Z++7wMc6I8PsWRT3uvwE8rFjxTkQSoSEFNEfnqzCPBZJJ+apEbrUcAu4ieQsP+ogP
hlhztTxFc2bgCpIQrNNllUJHxIV8VkgGO9FeWA5jjwR06A4O5qLSQabFF1rWKKNRwpDwP08b35o1
PPZzBsg3Dhz4eQbc/rDDboCbPL+dzvlUtvIj/3uYxZOhZXsehnd7tbVw6+RK2GGcNuIz3L/g5urt
XPsuSLxWXoUejzK0qxs3PU/36pMZUVBOdwpJY+6sQhiULsaqT/AQxTtbHxXKiQsEu3egFlrXqjVI
NXtADWADTngxyb9b97bdRRu+TnxH8JjAl1k9M4LvFXPUDq7knooG/0ozDLKRKsqGjFt1OnEA0z1m
WbWNv2KxcWXSPUvTrR/uoyWYWiX0H4tZGeEqCb2VO0HoMlzAfU/PM2L+YRO6cSpdQj5iG0JoHA0H
7VHBtWImPUIRCtWDRbZERH5t6p6U78Os9MbPuvDOqA4XT614VxPqYw5x3iOSGNVKLOpyBULdNaaQ
s4GbSMSv3S2hqB+bx+mXtWXY72wlD8SjxgMSIvETGBVV+mWmPbjsnVmmm5WAMF6GfPAXm0XTXL3Q
AoKItO9MZtT14ODHKqzDmbaB6lJqg5eOHCWZ2jXHaM9lP6TIAnM53PdbS7tGf3/ojz0dsyYmafiT
vKic9W4t0xVuEdt4iRhk4Tcia/XBoMZEm6xXBQ4CmuEf2Ps820AqHH/1ZJ5gqDn8B409EsNfSdpb
MQib0JMALExeLya275sb7Q9OHHOsj4cw+8ZdxthlFcdhzi57S2NXWv46R3+8Ko3gOXBAY6RglvY+
PeXwigGwlhR0eq3ZeJPBJaTSOaAFMC2zcZ2VMSNLCPAoYXml/WlTcrrBYLy+l3dWQeZs+2QeML0k
oSBd50OMU8ond2/VoLGZdFcUwJuDja/g/l62JtQ0jO/Vhe18JrptZx7YZmMqH8n/zTPIPbyPgTOT
eOrhbSDlnJW/Uz4VUR+ccHvhsujzFmEM/+GxUarUJ2QktGqHO8ULRLMBHZQqHNbzazCGgm03OyBe
/Nlvq5qhttDSWQAu3Uj0zeQwIHZd8JtQujeUeJCH7DWLWWgFQGeV2cjyruyzLAJW1XefJ4M8ThqR
82PhuCQVCzvG8qkwpIGBiU6P79z1kYUXVGbSVxXxeHkz7h7pwy68vSO9WYsyNDuKCqRFN95DKZlS
fGK5UmJkuw9KRsvm7Yhr15Iohg0YDwufaCSdmUcP571CLjYKYomKvIOee7Yubkyq28a3yIZ+Fm0g
9Wt8rWgKgEORn0CH8jbuajCWiJZ1PUy9tSgSuQANvCLynQgup5biWHrSIQzbqqX1dtvTG2kFHFju
CwdSjN0CyXMTQazI5qIWWeM0FxaIvLgRc0+z4fVjQVhKOGHvLFUMMlRkteBr1Zc9GZ6ZZXQwc3wc
UhOyutkGJI6wP1T6VoDMBsWT2dBJ3cII1g21Mz+8PzvAFR8khWxgv89kKz+RrPRPnLvca+kMest+
eVUvA5klViwuAMrDE9BUkc6FSV8FcexciJlLOYiLahw7WIdLIajMJQN30Mt2oVRI6MFYEOeHsD5x
BippW4GGK2j4QwN0SA8Yd27DArjijd8H5NaeJ31Gc5Q7apXTt9HHV8aUDNrzSRvS0U59eqFKcvMl
XAHTusi7VLqWFlD2hkqJmkT8wghdgLhoPWZ8nQRU40f9DpL3onXknmsfdO4KJ8s2aLeQoyMekgmg
r0luMtkuNr0WI7rq3Cox/Jb8Sf8JfYU+DX9xd63c3aqL555KIYDr02xDOYSc5VV0dfkDx8rENtzD
C/oq1KVT+e7oyVrzsNxLexAgmzrrRmkm0QZCkAoqyYFj0QEJ2bVDcSxDkVS8QNVTCUDXogH0xE8o
Nxytb5d04KWxASHjcC3Hr7kkWPiFq9HXCxdQIK4BTNHxZTXwHF2+oUjWD7JRStl1Xa1OOPcwNepL
XLvYTHIxNlPSHcMOlrJdhDovA/WFUpoAsjKJamqYbc8TjTAQTr5Gk+Q/llZs/Wzk0cAE+GAKuBZG
kkXQHQrleeg6AN4+oTjQge13uoprR0dELlx8w8yWiOoQ0gJVYdw31gbBmR9fWq5mA6JxSMsUiFt9
h/gxGD5TAMlU9W+ARAyu1/3z26NTqJl5rxi+wXlkCIhDWRldOT2Jw7FKKkWok2AtPXvPGZeXXYbL
4U8CHosxGJHc6fKZnLC1gzeUtKBvTi2JilgM7riFK4VWJwpY7eJ5km1pArh4dBbB7ETjgouCcx6q
MOM7AMT5N4thJUrJn2syKbKitj3Du4Wg+ZLSwajXgjJDJNqmaKm6XPgAAuypRLKq2GH1yp+XjdQ+
yq1H8hBnCqJqTef2lhVDmDVE7Axm0V2IipFwwCn5nyeSdNVvusnle2l5ACrm2x978gL9mi9czu22
cNRBnk9vLRKBDUwqQO2rLt2927C84CW/Jsd8seiNJI3pIriBWTSkIUFTREWy1yeckfxlc2kVbM83
yXifolavDWHbNvlUtMKE3Nln3iklPFAv7zfc30xxrJO86O+YY2wLSyyLODu8UdN8ZCCFsYj0LTSA
Y1GmAgUUg4OeodRsWBU/5dXGELip7jW871Bioc6K+xRk2IxBqRMWClOYqXG/dL4nEn2vTUxW7suK
tn/wVNJ9k42Yjd//fK4PdMgHwenxJmfpxOseerkGtg6d5UQ8JWwmaVMavSjusl4E5y+rWtS/LVS4
bGBWWgeP3iIzfqQ017f8LXErPWR5JxNes8JnSDSG8Waef37ot3ID75MO+Fc7o0YHMc7a2MXbGCaN
FFuKkVzcesWmhzV6fH0B3dHiTuiGcbatUYSKGq1+vt0o89ANSNjwcFwCqjsCYBo7ATQUamVwB1SF
GWb38RvwSUUGznOF8OO8N8Mvt4yEOi9r+PQMVyfHfC+xN/t4f9iaWy9k7A10oxPIrz9maDs46IgE
WAmYZW6VL6InJv/826T/8ovQzEYqh4C0Dl1d25Y+CYovRkyrAd2VjJa5SOCgvWQCaJ7zCXt8IYcR
moW0QLvjHbG/HM1WsbrOhljU6FJTPjohYK8k/b77W7UpF7yCmKHw1+L2
`pragma protect end_protected
