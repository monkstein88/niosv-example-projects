��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��~�"Sy�Fn���oL_�/~k�%�/�/:�ײ2�|PO2w�7Z�VƀЧ��^?c��fP��nԚq�
l*,�LZ��r]±��3f
%.} GJx� ���������ar�5�F�]�����)���KѲqH�]v�6?^v����r#4����v�]�52�/�u�t.���`?uP�J��i���vx����{=l�u�	ւL����(�f�|B\�	I'wL�h�/n�2�˅=�9�a�ۖ�0�~�<��P��4d�[چ��1�ݚ�dz�U��҉p�kG�\#���-���o�@��	ɬdBc^>�� -�y��%������h,A4��|�9.Ϲ������$����V*���\�i���+9�*8���Wlpo�/���v�K?�j.�·�5WK�\<č�������Mŵ@-��$.UPV]� S뾶��)����im�.�־Ek��H@�E��B�����e�"���������$�+��)�Oe�R�:Wh��3��Wa3ѕAB���'��)Gg G;���SY�S̈́�̗x�K^������'6��\a�9�J�Y- ��c�Eo���2S,�/ȿwh�|�&�{�);�:v���P�#?H'���/<���%46��*Ⅿ�A�,�m»�Ė�g���	W11�3t{$�e�qLR�4����v���غ�Gue'��f2�#.*��>F*_�c$Er��vUd7c{.Y���5��I��0ɿB�[��j8�D<�X���m/���H�q�3+ܲ�u���d��\��7���W���s�n���ԣ4mm>X��&L�z���F8��ׯ ���X��&?��U�����(���\'�Ia&��f�Z�8a��|3��'�d���0��14��gB7��yu�iE}�:TNZ�j�?�n�Ln�����,���~g �V]V����TM��V�
LP�_�#`�v��.���
B�k�S��g_��p5����nH}�ZLݡ�_#z{{�k�5@����h<�< �M�G�Mg�8ŉ�>٨(�`�B���{�b�~���]E�dOI��BpR����F�/[I���$o��y5��+�Ls�N�|3|�1�W1J1��c)�c��hq�K��uq�e�?�ErLh��-���*�r0�_��������њ�@KO1��� =�����(X]���v��� I�2�j��T�q��E��92��x]#��J$��iL��~�$a�2� 樖zD8(	X�����!�v��I�2�=�`1��4c�=e��i��f�C0uN��Ϧ�9�e��4u:g׽��%��\��J3K�=��`[��*�{!�j�;����#J��ҋ�O'm�� �m�r^�Lc �(��%�cw�#�6�XC,��P<�E}[M��3�kLE�|�@�dz[ər��ڼ2���N���L�/�V�ʥ�5�1aŽfv�.��|T��ȝby����ji�w��P�H`5C��5U�' ��񢣚�me�lD���G�hLQ�����ӓHH
Tq�ƵƯE07 �\8�����U���P���j:�� M�!DR�UÁ�|�/�s^�?5ӱ�1� ݖ\�D�;&e}g܅�}l>R���<�Qn�8����q� l���,t���)	_U	��Mh!ЁULA=l��߁,jQ
ɕ�E���b[$�o���1�٤�c�6Y'�1�uR�.������cCG���+��^�]�pd��T����{�<&�C��z$2��7_̃aC�D˖��D��Nj4�d6�U�	���Kx�Y�s�ʄF�X����񐞙H�/ t@M9X�a�����D�j�z�͒���V��M"�&5-��6�������ʿ_(�:�2�LG�Ա���&~�m+�jv���!]���ON(�$�Hh��Z`�g� �,2��ׅ �/�ų�v�^���}�װfدܴ:�J��U;G�P.�a���5�/��W*+¦�2��{^������M"���߃ς���ٍ��t��[�q�i6�mb���+B�^����,&��5*i
S�7��vGo�@/��zs��yn]�R�b�G�\A�;����Ly�֚����(���B8� P��fBtU$;�� ��Ե��
D,�am �x�J��x�{��ю���O�8���O%m	�1�kj�G�+>#���;Z�hx���g�{��n9����=X��H�Q����[f�AYP��0�U���&|�R�N��:n���ল�!fֲ2�ln���ڈV!!�&�e�h�J~�O�aax��$2�\`�����?A��Dvf�&��^g��E������o��(�	�`�sR`�CV�c[��/����̸���>7KG
]<��>7���8�C5�׼,�����=�]���%E�EӘ��8�!�)�'�4a[�7>r�4����uӳ�#yP.P�HE�32�j��9�@�X��o��RǴ$:��&�2[� ��~����v�O��{�6v�.�f���g}��?�i�;V�G�)(�}l���_���*�4�{:��V:n}��\���oG֣��hn8�Y`E���7��K�ZY:bv�z��>�?�[���5U�5uq�_���,*�lg����vuK��n��E������k���Hۛ����Z�9	���,:.�D�L�MDl?F~�1Ś��~ODG�·۴����^�D�T�H��U��U���|8x�vY�/=0u1�8�M�,J"o�����_�@:RſY�
56FB�]��B:e\?;	:�K�K߳N��":����+�%���2�w����ZB�5��$�p�J,��
u���/M^\�p ļ�:�`��al�Q�!�)е�����<�ĨM�KZ���&�4�n[�����0%�vO*t t�W~N���a����F�Ǘ�I!M�_'<X����>�
+��)[�0u��.�&AEH�oQ�r�⋜g����aS�-ia-�*��籹�}��<��69�������KO���b1���P^k��>q�U!!(Y����G!�B/��.J�3N�?"Ƅ���N�U�LDf?���/������Q;��R{t+R��bl��0�|���q�;D^%�����g� z<V
��`��H�z9M<�;�wj6���;M�qF�c�gr\��cO��H��.�,����JՒ{�D��^�Yi���=P,��n�K�;B�ϫ:��<7����0]�ru;w+�č��em�-��{T�,�(!e�\+�E{Q��?��K�I}<ҁa�ܹ뫽�4��:tb�����U�z��)ג��&Q���^�*}��Cymx���"��%LP�㰞eRaܿ���3<���^�#�~S���[�76W4ۿ�陊�γS6њגn,Y_@s�֋�e!���`�$�%�� ���,�q��@�?�V���+j�a4x7�85T{���r��������Q�Rw�Xv`��~��_]�q��r�=	���"R��c<�Ŧ�]ko?�l1���Y�ǂ�	����(y~��D^=o�M����6u�E���a�Ǘ8Ր+���h�>�f�Nd��S�"�"�n���N>�G�倯��|�]��󬴩�I<f��V�!��>yz�@VI%��es�5-�P���������B:��E!���N�cAH�v?'�D3Kq+U�� �PD`,���S�~��F��v��$ݹD�����1#2���a�R0���?`�����ou�m.� �O���[R�FtD#z��}��&�`J�����xa6��0�����4	���P����Rx�{W9�`	�� j~�1�3+���	X�*��'�Nv��ؖW줺EP���9/��#�԰�Ɔ�~�m��~��m�ت�"#{������@[�"���x��� ,��t�t�)�a$�pѡCUd�8�߀yC}δ`��iF�$�O��#~�o�:�0�M�V� !�62�G��{F���z��3�/��8Vw������c�@�F���9x^l����sq�tu��T�����v����:rYYCf��!(i�Bq�9i���u�D3���;t��bc����ڌ;R��=A� H^WH>f�ݳ}�������jb���!���#E��:�Y33��UB@�A�%7�38˚E�ٵbX����\�o�0x���������$Aw�8Q�X�-�W� ����A����̚6	�R��.��� '�MS*N+�N%�% �@�pH:Jf�wk!ZV-`CWf�\��4	-����������F�*��2�L��q��Yf ``�籬�0�����1�>�y��(���e�*!�gK飉At�$/��f8n�!�9��99U'�X�&W�_��+i%�?�r�L��jl����:$H5����U��T2X#h����OJT�	~�o�C�ټ�_��=��"dY��[�.6$$5ֻx�R�z��J$y�'��Ņr�ȴ���/#�i�|N4�+XAA狘P���xL�)�����Y�T�"�X8k|��>gaHKܐ\G����?�8�F����������L ��W/�0�Q��ƺ�
r��:�4"q�*�߱BuJ6��M��Q��Y���-h����I�7
fw���� G.��k�S�T������l������د^�y'r̒X7Fo����M��Ѡ��Q��,I��i����zº����Qّ)�Ԫ�����H���0dB%K�X��h.��J�>���5��9�l1��O䠳�RD���K��rƏ#�hп�-L��ƶYg ��^���P���DB�z�8r����&�/�P��=���3Q�zlwS�"\1{KS|{ܰo�Ę�/���~N5�.�$�1�o��T%Fb�m����K��_��Y蛶���NU�A�*��凱�ƈ��%��5 
��3�Hf��ل�w�IZ�k8���f���Y��ј�����ߋ�\@���1B������@�[��yv���l0j�����������ݜ��9!8�SM1��wtgb���ZA�}��7��{Mx�C�ckMۼ��c�E������vƹ ��mU��R�q=.���dP��KH��k��@Ɲ�����%�3�*ǡ����Aݏ�̧���Ӯ�ٗ�`:F��l�a�����%/�]~QsN(�Yy0,�{u�l̕�oY��)�^�=�a�� ��M�}���k���yH]�aM }ˠ�7����?��/L2}�	L��>p�Ź�	6��K���%s��K�Yn��Z�=Z�O�Q=�N��CxQ#>�F(��A�{��� ���w���ң��!�-��'�%>�87�C��{��A.VG��L磲���r=a�>أ���*�o+ˌ���-r0��A{|i�v��s���?�ա�P�q��ā �IbKӰ�	���N���)W&J���g���*���70�4�E��+�����&�`=+�j�g��O�M_N��D2I6�D���^��[�v�^��yb�n�E��e���=������,j��=��YT�B�'����~�ڭX��9�L+Y�X э�(��*k>��i�w�\��ʼj��Qp�B����._i��f���>�yV;��tC?�J$�Ci+��:��">�(C�X��W�n9irRw�TD��oh@̡�6�Kc9%S�g������� ���S![W���Z��}����7J7!$��(qw�_�tm�b]w?(t:�F�̴K�E*�r��r���˱��aV�r�$�Pӛ�[y>�`$�qQ�;DaE/"�nkwbuwO��o,�@{fb����.'��K�5��3��aD�u�q�E1������{[��>J�W�dx�p.�u���!H@liS�8�e�<�|����N�̾�������������rP>f﫛T�}��z��o$|Q�fa��G�+WF����DyAH-�����e*��O����*᠜mG6��me"�m/�ZW��=�/�oi|��8���7
�8\/� �U+9#w)K�H0�>KR`$�O<���Ȉ�~�|d�	���/R�؇?T|I�=����9%W�(�{+�d��'�e*ʯTQ~�Q��6%L����د��愨�R�su)W�����	{�>�j�Ư���N2�T�g��VB��e2�_����I�䱳��a��WѰ����{s�k��ݑBO�C�4�=��>C���z��ף�)L5��@V�������s��Lf\D������$�oq���p���H��HO������MQ?+Y��P1F]��� f^q	fA����O�2�yy��oV�\���F|�w��Y�(x&~`����|���bE�FD{
?��w%��	�w}/���#͡z�,NC�<	�柞z�%5r���]�-��c^m��7/�Na&+���������gq� -���QUރr�Ö�d���a�)p�dd1 3�|���I���=���Z�*��C�BL]ԢM �PF��$�AH���C_�.D&�^;�Wj�Fh�vN�[O�껻���W�-�֜r�^��ۏi����qL�0@o���� a���ݷe��>ݹ���j��X�	��V�,��v]�c�˷�=��.*H���}"��,c ]�:�6E����X�)|�7���踝����٘DÊ�A`4�)��kZ��U\�}�t �k�z�h9K��aK��I=��4_i��GT%&�-�"l�LT�;$���{�[�"���1�4u�B��O��ӻ�M�k���"��h�QTC���ݧ����0B<g�����<"��P�,5+�^�z�l:ci%?{ͼ�n�܍���N�0h$�� ݎ�ID2��k��9 +<�zۻ7�t�BwK:)u�E�yt�Tu�9��%wSo[$kU�;�*�۲ �
d�6*�C6�L��E�Df9�Y��wȄ3�X΀i�E��;׋q�������5FB���*"�Y
��$�0*���ԙչ���΂�4z���Ie��yUd���{Є��@�PJ�-E���P���!2�$or���5����Q(�^-R&�B�IIℹ��ߦ��饑�Y`�-��s^�A��M�z/��Ü2<�03S�����p�$�N:O�Vx�:��/���]?Ye���B
�vem�v�K)�� rB�����,��W姻[/%�2�����˚�Q�V����R�m��wtŉ+� Q��X��� �~v�xN:m	9`6f�P��Q�T�*����{1]��5(��le��N��܈l�Z�/�����[�A�enh ]�r֦=Z$%����� w�ِi2�����N�I�1ϗ�J��Ҵ��U�l��7݇��F��P��Wg�qNvF/�d2��0�7
�.���LO��v��ŤdV��Zx^��g������1f���ދ�k(�
��P�th��a�^i�c�O��ah	fq\��Up��P�z��	�Gi@:(f�@���GH3�۞�:������4dK�y��'���)\L��j���w�n������u!��ޛZ�K��Db�8.�t �u�R��vi�E��)eV��Ւ��d��p�"F;Oe�p�Ñ#j����yG+�Z��T�2H�����KP�^ֶ�&M�"���h����'�CHީ����g���d³d�^�������k�|�Ga���x�X~�,\>w�-�����>Eʃ�ۡ����/���! ��3���/����Kyu����Q�"��T$��?#��>�!�a�IE������5�`jAif���]B��V��wҋ?o"�VԃJ􆠥:�]��ŉ]�Y�a?;�����,^`m-Շ S��9%)�E���Nw�gbFp+7S=�G�"�A�'P��������1�����Qݓ&?�̹+
g�+~�0�
���~����p�����́����e��?뒡�Q&�Q���iʭ=^�����,W�B�.�ש�F�Z(����<#'��<k���;#4��AA�HG7�I�n݅�M����0��,�^bO���9��队���c.���h����m�
h�h������٢���D뤅ɛȁ7C��\��m$R�2�U|h�:��δ��*�+�����@<r�F{4M�� �z�G8p�]���]1*"sǲS�q�� 8!��0z�ߜ����ۃ��p�)��@U�R�dl�c��������^�;���1u�W��N_��9v�5�/-3���
��T��.R{"	�+溶�=�ݘ�m�����RIe:{�r�Ɉ�*rX+�������Y�]]�p����>l��	Y�UO�9���G����}�Yg~R ���?$e�Bd�.�R=��h|ܱ��)���x5VȲ�R��3�ؔ+_�hp�U����C��C9�S�[�6�F��dmo@�> �y#�O���!��'O���"��I2��q�"����]ت-�����/q|�?����L�1�|�dd~Ф�;��LΟ�.A�!\�����N���Q��O�UG�î��1PG���]6G���^{X,.��{uRJ;.4xBP�&V��3�@Ny�v��V;!�f!�� ��>pRՋۺگyK�F�QI�N �g��VЛ_o�'~j��G.���)��h5G�h�s��$�d�mQ��UssN�fd��rV�E��9�Ւ(IJ�����<L����=������^u�����?�v��HZ��!/=]ԣ�ņ/��ԸC��xd���;�|�̫�����C{Şt��SZ^���Z����Be`v8>{ҝ	�S�kowK�.��b��r��"��+@̥il�<z��3�QwR���5���Σ{7a�'�"���>�[�� j�x�0E�QO�����Xt&���\���c�CG�a�:�q �u���CW�@�KP#��]�|���S��y�q����ƾ�RCB^�t���\8saE�������dTx�]������G"r0M	���ʫ�F��?�!���h�B0y�"!|yj����JZ��Y�B�[�8A�P�9����}~�Gy.Aŵb�C��3��Ҕ����ˢ`ߓ?Tk-�˄�����!$��>�ܾY�9^��`nqO_�qgXr)ԮK(k)x��Ah�1`R���7Dϵ%��������~sU�����6�}-�׼qe�"����)ӆ� j0����r�wMΛ��g�C.נ1O�s?�s�OrY> ��\X��l~t欓��+/�� ���OW�[ED��� P ��r��b���F4��ZQo>�595��@ڞuZi�)�۽xc���{Tl��W�VE5����A��- tN�ώ0|�{$6����u&�_:���J�p�H�<�:���}�8��W�q�w�=��l���d��Uէ�i2+?+�o.�e1��Ǆ"BxB��4�&�hܐT^�`��	��zÎ���B���Ŧ��0%Fl~;o��v���<������)R��Y�!��;U�p̘%�Z�2���Z����I����!�ˋ6�9�y����������b��m��6`�G0�ּ��x�����U�c�K��*�2����6�	w����x�N0���$�����'��'VE���u�VĘj��z����>l�,'�u^�}�J����ls9a빣Â�� �q3� ����k8���O�J����Wb��h�U+�N{v��� ��o���\���/)K�>�����ϽV6�Xǐ��)��:mo�#����Y/Q�Ҁ,�~H�f;�~� ���Sٯ���aC�s���h��{Nz���>�>�/	1��Ʌ�Ք�[�M �U�m0%������P���4���7Hз<%�wԛֱ������j�<�!�6�&E`�\��̾߱�EQ�3�J�"'Z:!�5ɓ���0�x�/hQ_�\G�8�$Ar4�C6��ƛ��m�`=�Amn\m6���6~�q*:�)n�|�Z��v����`�r$O�?��UV^�M
�����G"ԁ��Q��m�G�}](���[�ٟ8t�X}<�.���?�(]�&G_�� �b8� yᔘȢ�C%���an�M���-��;�
~��P����;���Űw[]j�1�c�T���<?ţ�T�BZ����ez�P��2ʳ/\͏�:�1�a����`|p�)�YksT�$z�A�;�Z���}�:�S3������7�_^�V�E����p�zb����T�,������A��٤�l�y7`{e0Ɔ^����Z���s��:�����,cלLN��$�-8�4��Q�ݔԶB+;j��L<�R8R�O��4׉W����9�@K�:���=�?�m�/7�+u�e�_�{�ƵN������V�:��n���?��M�1x�ф�=�j+�A��0C
�9�O8�h�Ǌ��گCl��  �@yW},R���T����4 ��W�lR��)�A��O��ˣ5��hn���������~����x�*��� ��/� j�,�ƶ!����<�V���)~��P˘���H3�5@������Luk��Ќ�)Z�)������n�I7W���75��-Рk�H���㣩���;�rjJ/��ĥ����7]�X������ul�y��9���|a1�#��h��AKX�.����N��Q%����_B�?�k��\`,p�� �W�Z!B�tz&ė��:��uC�>D�&��i`����j6`<TI�=�n�T��ˎ�	�ےV�.?�sq�_2��/0�G P����"c����0��Yy�����N�?��(GiQt�R���f�T^�̤l' ��I3�_�Aau�޼�*���5%MW��Ǧ�lƥzU��E��[uί�,�G�ƶP�R,�n}>�Nr,�
�K���+�_[��sȜ%�ߟT�t��1(��~��e�:��V��Uo���t��6�
t/�rK�Jq9!��V��HC�����	��׏��5�,k��jri�\)!� �;8�����sG��:�F���N���n�������m��o��n!<���"�О;�5M�fH�C�o6���`�[4É%F<�uXԐ<k��W�v�G��#|�B
��z�p���ֽ��N���@#Sf����7��@q��y/�3d�e�GK�
Em�'���\V!

��q2�Jnw;�*���N�n��)p�#-( +��9͕67!i��b�i]���\;�t���H@�F|u�js�:��[o"Q���L�U�ͤ�=q'Qq;E%�+�"U#{ǅ�tg�>rM2��4�*�c�o��VSx���y"�^���W*�VS��}:^��7K,ʚ��5*FY�z!��o@�{s��y���A�a����}�L�Pђ�c���(��֓��M
�Q焘�|�l)��v5����~@<`��!�Qh������`���Dܗ)���$��/�Ai��Z=|O�xѯ��x$��yزi�s� �3綁��[�ѥ��iJ�6T|]����W��n�����i�'���g ��<��4C-:�.4i�Ʉ���>��IOS����]�vN4^m�2ڠ�A>}��Ji�CŗG���πL��2��^�}Cz�R\1��0⓰�P�9�@�����6ږ�i'���ӱ��^�	
���e��Ei(P
�-�1��`7��9�`�>��c�O��$�#T=>mȠ1����6VǞ��q	�0 ¾�o�l5�����M���~�#�j�[{�~��N�ۭ*V����I�>�xl.��t5:��-�7�Z�d��k�;3V��kP\�(�x\�9[-��N��QT����X��d`	��^�b>�vM���땈fR�G	zt�}�С�e��qoI'(��"�-=X&���W���S��`������_x�_�� k�e�檀�%Ά.�ɂm� �y�#v`��JOj� ��{��k���Sj�>8�ıe����@X��4�p��v��H�W��񵝉w�!*5Q\�U[<�����t�~�Qn��(0��T1?�:��|�d�ƛ�������W3�CG3����sGI2��`kx%����nUoJ�А>1��u ��_��4y������eZ=���<�ɫT�>Gk#F]�߀�ˊ(o��)�A�Wߌ"���Z�w���k۩�z�t%�7J����6��2���\b���	Q*]1�0�r~�Ɛ,��u���}
����̋��e�Y!0�B�zY�����Pjr���$В���5�{��Ӷ�Z8�����MT���Ԋ�:�X�ʎ�-:�S	h�~T��/���L��a��ԙ�D�uO���>���d}hw�Z����vƼ)���VFө�ݽv���"��C@��Є5�4��{核�����<9'��	K;b�U�<�h�qk��X�X������Z��>| y� c��#[�̝�=V�s8 ;v�)r��G��I��@|tڰ�`�6+\���<��j����em�F��2�Z�~��Z�6C��` �"�~�*���;9�t�#Z�.I�Q�l��%{�f�Gm1����Ǿ����I�: �9����o�����n�a�ځR�悝uh�&|��J�+c�����_�,�0���`�؀m�~dl-*����CQ)M��m�V ��rW�:�2�@m���O�FF�0�}}����Z��_�i4�J��O�V<ꗘ���͒����� �#}��P���-�b<�m� \�A7�y��ӟ�Ι��1�����'U@5o}u��|�.�i��A��*B�J�癣�' 9�r_�h���\���2_|�<t��55˜�؂�z�^�S�SL�F���!=����p/y����-#ӹ3���{�VY�� չ|'҈j�0���8��zs�x��#�A�����v���:����z�L�h��i^�\L�D�m�NH���g��ˮ܈M׹�̛AqZ9�lZs��e9g˖SA�DL��UCi��#|j������gOCaD����Y]��1��S��9:��K�F��m��(K��8�f�+��������;�QV؟ԛ0Y S�f�#�KV�<H�q��KA-��&�!è� �׹l��뉛���+����.^�Ba�WVM'<���rk3��C%���A������k�K�qqH"[��-�C"-��"õ�h.�1L�0�is��cP��2Mt��o��hL���>�^]/�+ܗ<<�L3����#��$��)��l��Y,��<��
x��
v�q�����]`_+��D�	l;߀�,�X�tC5���?����èW"Q��>x��C!"�kO:f���G�*���HWaIG��	?�gU:�^�<[:+�<��,��B�M�-~����M0� �����.p
I��^�l0�b��k�xw�#[1���i>�8<���.�>��Q<�J0��h@a�^^�c��k�%��֨?�b F��;'k짆� [kB2TG_Vk�I?B�Lf�\�H4���M�B�K����GQc�R�q2��}h�9����8܍����?��S"+ۥ0
�x�f�'�l�<Ԇ ���h�*�[��#��Ճ4�M5�ROŽ����.{:��[ �X�#r�	1/ϕ�.H��#�r;Aui&DJh�nq`JS�9��뿭v�_���2t�c�sL)>�21���~��� ���9���{����i�ܡĝ�%D1rtt�0���K�'g�0���s�������A�Y���@�]���h.��}���A�	�@��w� m��G�[p5��ܘ�d�,�Z�<�q�ʒ��f	;#�XV��լ��P0'��-�H� I��q-�q�9��g{�=���yv���^w�wG��(�������A��̢H&���"��f�^jI�,S��a�;E�͓bީ�?f5�˖�<���"Ueu�l� MK���R��ɺT%WLtd�B�S�[Є9SF��S�sy�֌�W)rFE��_��*H��@�n��e^�!���[�_ � "{9<�EYB�|L;vK�βx�^�]-N���1c|�OWeK��Spm&cWZ�

��g�0��r���e�R���/\���$�A�3�����u��"�@�G�᪐�Nq�V`}�i���a���3��&�0��*�QρDe����"m�*}��䲥�j��nL�p�=ZidP"��L�BH+���������e���,Æ[�:Os�-?s.=���}/��@�+�ր�~-G�% ���AZ��,�5��Ů\`��__�%�18���q��!5�Y+����V���	�[&S������04kTj&�f�Ϥ�ধ%�}���F�nQM<p��Gj�<� 
gk�"[I���r<>�B�>P_��/1$���#g��*W��h�Л/X\��k]�:��֬�e@M
��H�x[�����@ �ϋ��U~�m�}0FS`j{ގD���>�CX*(u�i���;Vc�G��V���W/��M��*��[8.�������o�ڋ��Ju�$���0D�8�@|��lN�~gV�аBY���6B7����8���<~�kM��W���z�c��1�$��Sw�4��ʪb���������*��V"�W�_��7�-�g��n1nq~^B`�Ē����2i��3���%��c��RuFhz~{xuv��Vb!�ED����	�O ��~��Y���X��9`�ݚ�uj���O�*6�/�r135��quql���?����b�����Nڟ��A��3��F���zs�3������;!�[��/�q}C���yh_V:�ê^����X��Uљ[_��O�������X�ߓ��D�z�j.��(���['��᰹xϫ���+�+O��
�a�˷V��f*t�r��M:��:�Y�k�c��B�t��sG硝�����M��:m�2(�������38������n�f��O��}k`�_՚��xon;~㛕��(i�� ���r�tܠZ��-*y��UU���FP���sy��*|"��'Q��ɰ�C��D��?�F����C7�.���(=s=�����~��jM���̪
A�j���5gj]0��!Բ��խZ����S^1|�#Ed�9W~�,I��;p���po�5��ݣTRP�-n�z���	D!�.�>��em}��}����g^W������p�x��<��#�����(<���7�C��$n�lM
"+����� ����qi�'(Y4Mݾ�
R��h������rc���ħO6U�x%����\��<�a� �����FQ2׬�+[���-��](��$����)��n�D[���'�4q�#Ha6}`�Z��}	�,�T����Y(�If�Ŷ!T��>��w�/X#f{�%IN�x�1] �)ԥQ�6��dT8(Җs���D��R�5�8��e��*?X�/=` Y�v���u�Z	[���Q&�l̻�	�1@�ַ@�I͙0E�0��L��Z��FYi�/W��'�����,��q��;�C�7RǼ�:�=�$g���d�dnɂ��x�@cw��U�i�i_���uv"�ȍ�m�{��3+�����!����3��Ò��F��գ��r�'�J[��f]�vC��6����F��n�"��[�Μw���m��QUHݑy�o|3<y<����wB�`��u�/��A,�e�0y�����d���p�ʑ�61�KN��{Kn���D�?��ޜ���\D�KqXW5���ܪ6��}�>�4�f�,�쫮L�3uW0�`�O��K�K���w�������+�9��W��!�8νzUN_���[^,F歃Q�L�h��^��k��f��}%��$�16�@��7ݍXm���jC�d�	 � �(CX��#һS
��S�!,��ޯ�C�
�z�}/�d��U%5;�H���|P3�d�f	���X%�Z��ZwxF[����#�E=-���V��ne��[(G�x��f�'�>��v��	���=���k��<��eĪn�� ��s�ɏw�~:�D��Ф~l{����k���9x<�-�!�<�T�өѢǛk������W%�|V�D�4���ҍw	6�/Z�I��O̱~{߄��=�f���oW	,�����0��j�#�9Q�|ѕN�T�o�[�
$�7�9��7���҃j6Q\� ��9I|7�d�(��l� �5�[�h���CIuIM��O���%�~!���Ŷ���U}A5���Wl���V&ۧ�R!6s&��_1c�c=�������x���2����#��$C�.�@~�G��/���tX��i��$ÏM�dc�;��F%"U63؀r�l���낟2�H[��M��
MTV|�����a���Ӣ���ݹ�����<N<r�=�8�.CP�ޡLL�����c>tcD�o��F��.��	�Z*���pK�K+i�ԉ�?�^Tb��(_���d�4��ᕑU7$ȵ�� W��Rß9�?9�;
 bH˝�|B�C"��դw�G@H܈p�t�!�|��l!�����e�
G�׸"��������f�$V���]p���-�q�;�ݜE�P�,���w���Տ�Xl���A�p���}
mY�jደ�%9s}��ZY��|i�f̽��֊,����_@3&�a���3\�����΂`���Z��0G>����Ϋ����G?3�i��A��%2>R?�?���?!9:�Ѓi�\"��4�[UԆ�o*�J˱`	,�6 �,���D0�j�@���|F"�%G���5�ΊI���4+:T�)����|H��Z�sx�5��`��eE���g�*`�H���4tE�|�Z�Gq��HǊ��F�p|���aGW�R0wڄ�����*ݒ
�h�.�2
�ܭ�f̡��|����p��AKW*����g � R3g*�"}���ԇr'�!1�;�Ok0���b��D���l|�3+&M�F��1��b,�8��
�y�a�����#��}����[x��A�e��C�j���`1E`�sx�,1���IZLҬ0!v<���S�~0]w�}��=���Ħ�6��R��W�7�R���R�ߦ`ԓ� $ZWw�Oo����쌑>/���}�*�0c����P��g��~k�:c���+>�������o���V�O�&�1-��b?��+�Qe�(�(�-Ӳ9�B:烥g�)��7V eοkB.W�jY�X�m�BP|�lD)ZB�9=Eݤ��4J,����{H5-�3��e����e%z���	,q[����?�W�Ԑy�[��+��`��UۈU���N#d!�	�+��0�$;m����Z��3�|��·��s���"2y��ϥ��%���Z[61��ЛB.�\���6���k��/��/�7�z�C�$��q�4�f�˙����u���}2|Vs�+�Ю>Ѯ�OI���&�c,E���	]$�#�[h��W��g����=|�mw;lIk`W�^��mrD�?>�1ؤ�,�	���@|>1^�8�,�TJM	kN��Xz��MJ�+5���g�ߗt�JL�Ac�L����y�
;���#�/�
����#B��-֟�驳iM�v"�V[ɫ[{ϘGѽ����4��x��%`���:^�zV���j��	I�b�wV�>�&�)�E��K3y8�&ɯ��x �X+N����7�'�ϗ5V��VC�a\ȆU�����m�����2��(��mY5��	IA;��U�������`Q6�E�����"6E�`���%e/�.C�;��ޞd��y_�A�c弃u�o�������B�:	��%���\'���<��RO�x��N�fm������
��B�����Y��iX�3e�+�w";�(�'	g��=��u�&����K1��藓�d,OMѹh���^���Y�Ű���W5ȯ�r^sB6��7ڼ�y��Ć�Я�:�ƒ���O#�4���"�2sFM�*�g�*m�:�yIF[�v6�,��l�A՝aY�S~���,z8�p㘧�5�D}���ݕhz�*����3<���}=SV��|�C��8)�R�Ơӆ�K7l5ww%��Z� ��|^>���;���L	�������\�ib��v�U)ϛ^-��J|�&���� "�(���p����o����� ������u�n<����w)icuºx�k���
h+9�Z�T�� ⵣS{���m��������Uޏ71��4G8H:��M�[�阚����:)Ĳ�槙��'���� =&7dv�h=j)��3�c��u�E����-I�Ί�F"x��+��x�� ��mU�T� �c�{�J���F�:��<�3iD�9sZ�J�
:ˍ����w6���4������R謎�����;��T�KD"϶����m,л��w�z=u�s��C�-F�h�&a����n,�{��<�`Xz%�a���c��� c��n9<�Y�2��Wn=C�'�OFazی(>I�i�/>ea��*�(�N��v���p�ˇ��}z�@�-S&� ������Mey{�c̱��=�I�\����hK#҃�t������7X���x�䨽�K���?��T�d
�M3?]Vx��d�%���(��6r�<0�����&rd� Q��0��;���.Nw|�(���6���X{���$��� ���[r��2q$c����Fx���`[7���4-���11��rrX��@3�ѥ��jQ��N��_�Z����Uh�"��_�[�`e3��! .�%�	+��t�κ)n�{��>N4;���~!������+�G}-��F��l���BU>U"���-���!�� d]U�#ׇ�"��_�JW�j�����s���MgZxČ��J�#�>_��=XawSka��1���D}.˨l%�>�wS��62�~D�.ȾMΡ�lR�����C���Z�bwO:ڀ��n��We�>f������M���ɽx^�^.w�R%�9��KIQ��.v���:g���bRa\+��C=ϗ� ��?`�<f�0�u��z2�){�c�m�K�`ȑ���q-��|�����>&��ٖ�b���]�0��(����Ȏ��uт�����@2A���.�D�2�P�mF������b^���ժ�Ǝ�Q���`bA&Z���\z�ǲ-�"`�aH���@��~�}�(�-�y(��^Y�r���J��"��f�+��f{�Z�0�H�T�Ic\cp'�ň��ˢ���C���ƞf�ćZv��E1������fM\it����V
eD�wL�����$��^������}�N���S�n��!A+������dy�R�
�p�	TdL1�8�8�6�ʳ�G������N�����{��g�P��Ӂ߿����d��8w��T��VKx�JO���)��l�������'7��K�'���r��ɞ�Dj�]��8��;�E����������-\�Ž�F{ �;���rMc��5P7���7A<B  �

�	�cx�4����b��{2��"��<�b�$H-�r�t������3B�'($E�$��7���x/0ZBݥ�ed����Z��l��c����V����L������ A�����$ȅ��ɛ��7&~s"=.B��y<4qϧ-��3��آ'T+
��(���|y�sHL}���Ia�\Ҽ�����pҺ�`3@�
JL��+a'UW�}o�����JgT(�a���J)|�&�����ia�(Pʬ����k�׫�]P��{��Rb�[,}���r�k�p\�A��'f9 nv�.�D(��q������X�� )U�����.1K�x�oOٚ��Q���W�J
+����m�����)�V`U|��AkkEz�3x�y��� t]I�i�<�W��Z�����0�A;�=�������WJ�]��G����ۆ,7�α�I�ı�'�,h��Pp	&�Ì�[]�������;�}Y�����Th��.�R/0M���:m�P��a͜�J'n���^Qgs��y�K؀�<YV��\,��j@�Y���>��ӄ�z��{<�g���=?��ڧ!�
����B��'�������@3�M����Q��x]!+ڊ�R��,V4���6"��Z)8D	́��`qb�X�6[d�C��ĨG�#�m��: ŵۖeE��B/Nƪ��y{C�<_���8��8��+!&�Be��c�0U5��� �'�-�R�V�6�^>� ������e&��3B)�(Ƥ$g���p9ɐ5��l��	��㏭�\��A} �������/_�!�p�s��3W��=�^EW�Qm�u~c��̗��v��v�����?%uW�^���x���L�Y�Q�d��D�%+��b�}I�S��ؙ��VaU��F�om��~Ɲњ��a��7�s��p�5Z���Ieb�k��O�P��J&��˄��RݫPT�#Tɹ]\�g���4ժ�ח�����(T���Զm��<��C���6���qa�v��!��� ��J��dp���g����1�ؓ�������}�xL!�+ӏ��\�$P��Ȧ�r��M�Ϩk_u���h���Q�Q]�æl�# :��Cӫ�W�ͮ��/�ɇ�o��Տ`g��u��-(ga�+�/�n&���S�����l���t�4�âu*B�:
�{�AҊI��2��k$8�
 ��Ͼ�5��:d�u��~q}`NYη��ȱ�ѡw��¥̽��l{]���:�W#����|0\k��?+���xH�:�r��;��cf��̔���r�u�U���-W�OW��[j����W� .�2mJW��ۮ:s�-K��4���Z��� m)s.�+`G�k�Bm|�����y��X��pe*i:ӧn�֋ػ��]=�~��'��!'���Gd��m��;�=7 t�(�;�+=U���P(��� �{�=�F�Q��g{(,,�n+o"�p�N�1�wg
1��8�*�u�V閒�@ׄOK��'}(!=BΙq2����F�E��A�T'��u�-���j�?�� ����Dc�_�w��Ʀ�w/�d@=/[�G�W��+���T����w�r�j=0���8vX�;v!��?��R�w�pltى�ņ���s�X��^Q��k*\C� �T/D(PB�U�qh����Ho��9<�2(��.��f�q ���ۦ1]���П�u� ��N	�/*$�@�x�cF�I�-n{�*h��
xZ*�<�	���}L�hVo_�<Gbt^X�x�B^R��& Y��.N=k���}x�
_gi�LD�0�3%;�|������A�8�����_��СQ6���fĥD��#_�Ǔ���w]����]U��y���˩�xVw��=�(q��r�:�Q_�F�N/+�4,�F���X���q��ܓJ��C�xc���I ��?�Y���i�Zvt�<����Ul��P���r�D	ig�E�?.��MIr)�ڢ �!F����:�268!\�貪��dA4�������մA�7��S����n��P�Dz��ƖK����)ߋ���	JJE
"n�����Ƅ��6��}�ڕs�/x]i�(�4�E��t����#fb7���F@�Mk���(�����;� ���h�	. (G 
�mx�@����UO�-�8n���aU'�{)��9���]|YQ�y�WDe/�M�������] 2c��K��9Ձ�<.$$]��-��c��:�gE�LaVV�FX��b�D����~ kU���!�=�[�P����~�H�c<�F�����^��l�`������; ��HhX��օo�
q��L�w�� %X ��lgc�H��C���] �k��)F$!DUH�d��1�<�-Y�J%�%9a��d���
'�c#إ�|�� �1�0\���X�c����� S�`�����%���5 ��$�����kSZ"����;x+~�����մ�\.�����B%Lx颉�ػ���U2�Der�`�M��7���䌻�s���	9ٚ)�����hQ�Ж+�z���wI�^�?�2V��sV�ʵz���+GN#ERg�Y��*%vUS�BFx�T=��@l�f��P:-�+���u$ϧ�O��������(�5zHP��C
�����8�$?�$�4Z�E2U:ɂ̈�(>´z�2�a� Տ��d�k�]f�V��	R�;*#8�<����9��C�Σ��g*E������J ��{��G��\و������"=���ff�Cp��P>��5�0v�|-���K��K�&��0$����|���5���`9v�B�
p,�!�#�u|�-Ť���}�?<���S͜�6}�RF���ZL:���uq�=����9L)p�r��ŵ��sunf8���Җ;�Ɠ��Ï�H��ZQ���&��m�U�Pmd)��`�4hH�y�9�p���^e�.g�MWEL4�g�>�o�R��x��(��gL�4����U�+�$��z��Qn,����fbҼ��vm�2�a�V��%�5L����x����ǟ9��iԘ^�}_�m+���3֑A��P�Ψ>�ʑ��\��X U68����n��� �����K�xP#�DV�P���a���^��qQ-΅T�FO��	oX�>E��{T�9m�3�$�V�T���·���ߩ)��ob����1d�j�$!���[�9�3=r~�'QN��隓8l�#0}�	ฎ��^��[��ء���3�)t���#~s�ӵ�� �חm@m�0%X���[^\r�S��T�;K��~�*8���4#��NdOO�TmLߨ��&*L�\Ԅ%ɍ�Ћb���G��P	.0'�*��7�OW�z�a�<�:����n�eX�^��Kw��#� ��w%�x��p���F�ـ-��Zg ՇB_��3��5{P�&j&�,}��*�<Ie��`yѭeռH�rU���cL]��j�����n�_��^-Xs��>�N���1ATF����w��f/gw��xb�u{k02�Koq�K�J=��-��Ȃw2J觛��`|5��Fx��Z�����?i�"E��q�oj#�M��=[o�6�B���nyGi�Rk��g6��b��#���]���R��ݛ��'���P��F�ZKd|hYN���AW-��va���P�f
U6֝�yj*+��dhġ���,�=�o��xe<O�aO�ą�J�1�~�
:���h	qe�|�B���#��U+��(�0"��+��2Lf���RN>�Pht�m8��L��w⾱�&A�R[ʟ���W*���� �v��0�3:��&��h[F�8�hd���׀�����[����P�΍��	蘷\��+�{���z���\�mh��V�ѡ�-f�\@�X�x}����t+z-�	r-e���/ξM���3�P+I�R��6
�V��oi����5q�:%G]���%e	��'ih�t�U+[5y_l���S0�'u5?�ٿ�oΨ E�wL%-t��5l���Uū�ޖ�l�zH� �/�i��ۑ2(UrX�|�yױc�Y�~9�U�E�9ÝÆ�	P��D���{�(3]h�V�&�x_?���MD��� Fx~��7� �[����MD��L͔��"<0A��Zu.�#!�!�ı����'�"�!�,?W|r��߀4�& �aj��t��g�L�f��)�^7T]%�C�����w|:a��F��{�	J�9�~:�������8���@EŠA0MnǜZV�?O6�Mϒ{�;�b'k
�D��]�*�8NĘ�CN�m���Rܟ�To8,i�+��t\�_�1}��PE�Jl��[yľ[/�ҤR*�t�^�W{��LD���e.۪ߤ��THwdoq�{a���,D�����8�����ƃ���K�R�})��SR�bV��������Gm(<O_��T"��ی������Q���p�8Ҿj��i������Ú��Rq�]oz�d��+�R7��հ�x�]w��s�����MNs>Š�֊�.s-�q���W�[�إs���l�H�T�17.�o��+]�V���z��Μ4�Z��k�'� �7ٽ¿b)�ƚ�Ŕ�  'Y��U��W Ö��@�g���P�O`�J�O#�����.��yNb���H��v6����$��n�1���?�k�G��~K��?ԣt��/O�rr{����l��y�w]%�S�4"�<�n���iڼ�~���(]�2��T�s��ɼL:� �����R�S\"��l�+�?�i�v�jʲe��_�H��C���ݡ{z�P����)��x\g��7�M`=�s�ݛ%W����V!�I���A/*�#�?�#��������� ȥ1�&���Y�^Т�`����+B�>54gڛ��� 뼉PM���g��m6�^��=�G��
��~�pzK"��ذ$V�풕t.Piy�X�	�|ti:��JL�,�vJ�T��o������^�"j���F�}����@S9��p�x�����ܐ4��sh�
���� |�V��(�]���>��	P��"���+@]����R�+����5x @̯ ����!)OP��zzY�����P�{�|�X��˔Նd�g����y����G�|Z��1ary��W��^�����e���e�j
�7M�w�9ޥ��*/xz �V�	��8!g\�wz��n C��57�ƢL��aO�L6y���𠳫d�GYKHi����e�Y�i�-#}����\�SaCnH>�:9ץ���R��9#;�x��V������Ֆ�߬?=$)J5R^w}��?Sէ�sa.*�Ds��7��$B� ����0˴O8lF��#yJ���j*|^
�		�����	b�>�z�M,l� �=��Mm��Q�B3�Nw]�@<dp`M@Dk�q�3�Z-�1Đ�,���pM)��E� ���� {���!���HQ"��&x+�j�s��5{n��"� ��'w|[i5]��Vb�lLT�Ќ��a�s�AF�&��B� yd�n��,�Û�|��L���|+9(�%��� ����.o�V�tTäML���-̷��~�y�揣~@(F74qt���C+��/�b�������o$� DG��._׃ˉ-/�hN�a����)���M�Gr�Y
����=0!a��p[�O���W�����.fu ��/��p3h��O'������zCf��!Q��&R��	i��l��|�4�f�"���J��ůW��tTi�����3����n�znڬN_��@mʱ��0a"G�&�H��	0�^�z��$b���I?dc�m'��½���~i�36R����Kphc��G��!�Foe���[����5��5Irg�5�*t1�?|�����uu~�1{w�pN��M^�ܩ�	bwU��*3�~�`h� ����,�Sz�A�x5k��ì`>¦z0IF�� (Ѹ�2#i��t���R���F"M��0"܄PxO!��Fi<5
���;�ӡ����~�&$M�Â�Q��YW��?|�n��s�0�m�|G`y?г�N"�߁�]4��_�����/�1�K�I�}Gkw�z<��8�d>�F+k�<����b[��Ux��0�07�~�l�ʂ�qU����@��\�D�W�Ǟ�Y�����`��Eμ��&Y�Z����y�@A��fP6��2b��{$yd�~ӄ#8���D�Eef��0��Z���ޗ�v[�)���,-��O���HIpt�ֽ�²d"�> AXT����ǿ���`j�W{�Ej�P�b��q�/�0f(�U�X='��|%XL���b��@�|9\�};E~�_-A>���xL~���v=VH4N����~㘯g$��4/��eRXr��'��'-��쾮'�
�
�O
u�]�ܿ=`5>���5�n䵐��`���Uf�V��Ҕ9Ԃkf�J?�|n�ò� (\�k���������� ����V~��m+[%�ݛі�������A�a_3*0�*4L��9�g�V�e�Ɔ�}��a��&��a�(�8��)���И;:��~eٷ��5���cyi����4c:������WP�z�x0�+d�kH���oiHյ�|~�mm��߃^�Ϧ�!���W���~%�T'�ez���H�W��QA�KMd��
~&D���GE�i���A+�����*J� ��"��S�{_���;�^wVtd�M�R���U����g�$���3Km��sJ��֕k�!�}d +�� l�Q4��`6�R�D���K��J]���pR�A��{��%l�
��M��o��Tsa�
n�h�~�As�!A��7{39��;܋m��="�Lv�{"u�՜����}��OR��Z��J�K�a�l.�د3/o(,�^(�'��=?J9S7��^q�E�,ݥ���O~�6B�����"�g8 ;��A7k��1��3�%����}��[ɥB��߷�|�p;J��=|���[۞��ɦNCvC+w":�-Q�)�w>z�U��,;3�<F�q�|�"p!�t��yw���f�T��%�mG���)�Mi�
�;ԉ�Śc�(�.�s�/H/�.��������@��>�@�e�T�t�/�����VU�6�+Adr���	��4gB.�!20�2��ؤ"��dA@t�g���4�(���Ęch#?8mva@�>I��B���&��uu��N{W,;�ˣL1q���Q6ݏ ;İ�������0���z�Q��P#웡��X����+Q�,�k]%�OTg����m^�R�̒a���@~��W��u&�$��@'ןM�"ч)���4�������){�V��77��p$��$�zϽ������w=a�f�����l%���L����D

E�"Ƭ!t��^;�d?��e+[%�܁�uZ2d�C1����'�M�s/�В"w���h����L��P���A��RE��W�,eQi�����$p��E&�	}�3��f(}Ȱ�`=e��!������{�yä�ښ0MӞ��W���c6<��6ؠ���a��d<ib��s�(�Ӏ��⊻|s]d%�}%�2�V��F~G����;g�x�G�HrMWW4��ֶ�	��wF�N��(���qܰ����,�%��(����v�����"( u~���3�+��X���]4�-8VM5O�fxu[=k�|~)��̣�+r�RK*kL�K��x:pf���&{�^'O����=�HH�.MBR�w����FT�3����%��+H�n�Vf���(wj�֟���<�o�+�[�Kt�v�9Js]!�������&`?\��p����UNI�IR��jٖ*��ڄ�+��
�j�<�����b�f)�#���'��MRf9���`�7���wݚ���u`�/H�W��p:�8[4�f\4e�E����T���?h}��4�E� �c�#"��l�(��RHs����ʩ׺�����0|0��Ç�s�ej�$/��Ȝ)�2:�Mx�S�ٸ���j��O�?rEzU`Iu�м���Hj�݀N����b��8#�ʐ"sθэ ����^mZoeb襸����d?��Ӿ@��2ǉ�|���ob��2��IC�3Z�i�q���)��_���K��7��W8�#�P�x�\���'<��t�%�p�F��P����o�������رMG�"��Cc�v�}�;�OIs�,2$^V�f-�M��c+�ڏǲ�>��Qrx�16��Q/�F�Ņ�0H��oe�����q�	7]år3��wV��zZ�4���,A���],w�t�������q�L��������N�X�:z�H������+���0Ŗ�C�L��C�G`�t��;p��[Z�#�R5���
e
����df+_эm��Q%�������,�F?e��!����>xR�+QY.\�; �U&�I��I����e'�F�#ٞ���~	�&;�a��Xd�=F'ǻ��*w@��h,k���ހ�5��t����0�����Ā���7��~Q���vѪ�7��倁���4%;
Yo<���oh�r������NLmO�5��(+׌ �pc�V��t!�������V�ܸ�#��b�x㾢��7V	�g�`xrW��}��g�M�r��p�ִ�6��ڃ%j��ȯ�:Չ����@[ЁD�;���FU�@[h�;���M*���S�M��W�:���R�C�z�N�\�g�z��p��7�*���_��&�#j�R���<�;��� �N˲U����K��QD�H���}�>���¸��¥�m#�K|�BOwAB�0�
xg�P��o9�M ,��M�w>�6ٔ�M�������'��)�|�)4��h\e����=���ῡן�f2b�[~�߆�jF��b�?�-e�Ճն�2�.Z�
��Y-Xr�_S7f�+���|��h�.%��e"	��]O'׍�i����a� R&�~��f �C��x��1��
s���ŝ1�͞�B�
!#���x#���~Y�:�Dӣm'|�cͦJ+*�Ծ`;�%��;���p��c+9野���J?��r�T�cQX���i�� �ٱ���9�TS,��Y#)@�����&�
�7��o�9���QWU�E��?�o0�� �v*Tv�j�+}��Z�]��c��^����
���>W<GĎڻǖK���1�/yY#�?�bc#xj�ˤ���qd�H{��"F��7�)�����N��n��f�ǡ��TOB���N楗v骩K�Z2O��H� '"I�o����/�aU�0K���0��~: ��qOtL�S�Bm��x7n�_�շP9��$��/���d;im����Ħ�`�z� \+�t���;�5˴�Ń�� ��4�[��ɫ  �����80
A2�n�d]uQ�u�X�|�������$L��g?�N��4O�fTW
qiIU̇�ߨ�y���ɡ`i�ߠ=m���D�����D���'ʪ������%������$��'�`��v�([<�׀r��	��T<Ľv���Ev뷈ݩ�Hv6���fA�1��������^��=_;g�B�	�W��+A&t�#�7!�,����$~�k;hA@�*�}Rubu�g����T#F��8I���wgM���IQs��i�e�� �xb�0���K��q��/l��a���S����B%���3-���rO�$�u^�e̥3��Gl�u�$��T�74���5L�lK1$�@�ݗ���ZA��z��O��I�U�7�D�S��r�"�)8% �z�\��vqF�N���)elZ�VDw
��E��W���mJp��Yl��ioy�M�"�D'Rg��io�I.�Ê� �B[	��
oXJ���� >����J �더v�k1������3$��7ʱS�VK���Lu�0�TQ.�P�;I��h�/*�K$DtF�[�x�+j�qu6o"IV�7*��'�jJB�B,���j^�k��*���E����a2su���Პj������y̎���WlM6n�x �Z"62L�;���=�����:ϵ{H�.�B5�x��2��!]u�n�i��O �V�.�G�r����uQL��fzg� ��³��VB����	�ˤ���0��y�)�tI�l�1<���(��N�$�, �Z����˛.�-�&m�v�b�r�0��lnJ�������{*��v��V��·u ��c��`���Q���?�����G�B���Q�uDB�<��2�7��5�ZK �)Y��R���H���0��g�Ee�u] FݟE��g�L�e�Jm��v��G���DS�S�b��M1ƘTJF8��������me��m�#�����Z��G�~P7���OЍ��h�l$�	>Ȕ��׸�"'o��~ 3�0�0E��;��6#�*�O��?��HDx�|�N�L�:H=J�J��:���\/*��oc<pRR`�x6�?n�j�.���(��_Fz/|OFb`ҦP���^~�c���H
16/�2��R-l(6����*O�R����*�&*Y��~U�M0S�.A��`#�^{�S���}�{�xR~�Tc1S�
����"�$=������ʤ��Q4���n��'X��"�-Ȣ�-�(�K�-x���p�Hu�� �/?-g����~v�zD)��Qm��-(Td,��؈]֨��:`�\�`�b��&
����(5!�����s;��q+aS�h�W�Z)Ӓ�#�H���Ӥ���,�/�5i���^�	d��#�X�	�wn[8�"�GY�	 '��Y,�sa��!��a�we9j���#i\��3C@���+�tX��m�����?�؅}k���jw4�Jm0"n.���!�Rؐ�'����N6�XE�p�Ϻ
�h"D9o-T�	�[�����U�:5�k���Сs���=[0�H��<����hiե�4x徦U�|�C��t�����6�M��!�_��P�2HQ�ĭm�Y�ܧ���;�`&��(<�c
ݯ� �(�q����8��h���7?e:*R�ȟ���Pw�������dB���w���,��v�S+]g�a�����~�	ʤ�8HX].c��a+� CO�}?�[��v�>�_��[�K��(-j����%��A��s���t�L�ggBe<W�;�D�H�a�3�QF+ -�7܇�E����P��"�5/�Ÿ���8������r���ى�����-�4��NJ�3c��0Ԩ֡�T��-H 83�M�b�Ѧ=X۴��ҔX�Ro�%�������<x��p�#��0%L:����x[%I�0���ɧ�Q�0��7v�����e�Bp�`p�C(����	:�k5��,�)B�:�?jr�4-���29����v�V9xVf����Z�,US�
���n&�?���\���,�h���ւ]^N�>���qw�'擈��N*�*䗄V��46��2k>���+�\�b$�)Rp���	���u����8{�+S�϶�żGnɡ�޿�S��Y����P�C���r�p�X�I��P�Uh�7�U�8s�}Oxh�;<���҄������U)���L��ބѢ�鸐T��\��0��9/b�2�|�7�&��s)��+��:��hO�7Q�@�������[���E��+���=� �[�X{�T�^�6�)�y����hi=�!r�� 3�큄E}G�(_>Eє�p�.H���ᰲ�7ot�m^gǠ:u@�����1�������}�6VD{V�X����@��#S��s�b^i8���A��g�����:+<�O�K���kc�&�� ��������M�!f�\r�\�N1Q�>��b*���`��7�}��?�ɟzt�F��o���h��u��3����K�
�1����$SؗN�����!#�M�J�T3̕�v`�ftg����6�8L�U��yX�4�`����PmqF��;O�o\��>q�ƞ�4��nEz]t����k��-gm;	6}B?�0Â
U�~L�i� O6�m
� 0�����D%
Ռә�%U׍-�?V\c>mT�d��u�RE�)x7T�=�Iv?��I�E�˾A)���X'��o�\erP:zW�1�,��~࢓��_�L2C��t
ǭWw,s՞��L���r�r�>���ăS|4�����qu2�Ǜ�*4��������9�p��l�/����B�>h#ǤZ��}.��")s����hs�Z	�����y�!w�z��E�Dx:��s?���p��6�߬2˺k%��[��S��ٍ8��k�VtX3��Ł��?#C6:O��F�
x��9�L�3�A�(�}ai��@�-���z�q�^�g>�V{-�g�B%���Ƙ1�)�&�ϨK�����M��M�|��G=��t��y�h�&���N��v�Z�� i�D��擨,��G �`��>�/k'G����(��;��я��e��MgUY3J��MEp��/P%@1��<%[F �ͥdTU��Q�#j��eJ�(+Jp�^��\��](��T,u�
_�A���m��&M*_,��(�G���\��ţr��m�N��d����%�`o ���� �Q��/�`H� 
��]�%'Y�I���OF��\6
�hY�P�	W|�C��$=oe.[1	z�[���C���g�o��g�Ak
�v�����=u�-V���R�(�A��pGA���x�%���;�/3pk��C΋��Я���0u��Xs������0�̰�7��h�����K)Sc��sp�j*����8��x'�	�� )��%ϙ�v����6���J�1n����ϊ��j�K�5-M�#9��`�g��P�T.�KA]!h��Oڽy�!B���㼯�Yvv9��8Jd��R?����h�������yy�g�:�4�kLqh V�h�Ք���"�����|ǈţg��|w���pM+?�d�$V��?���k@&��~��[;����>Y��eX�8IG�Zc��Zջ�Y������b������k�����A���,O�����5oLI���䥜g	��¨�<B�RK-��p�\wZ9���.�}�g�T6��%I�l����D嚥k��@��W�=�l|O�U�YijnRp]�M���|P��t�}#��D1T0|��@��`.R�kq&�|��7�p�{�Hє4R�{�s�p	+�ÃZwm�L�UF��o�9�LFg�+�������j0D���I�����Ծ��B?:N��&��a��J?Q�J[�v���7g��Lݸ��6,ȐK0���ԭb�Z��Z�^�V�m��y�ު�n�!����Oq�A�
���|�5F�tn_@�Պ)U��,>�<$��=��J��(3���'�wg�~=_�/�$�����l�����ͱ���5?*��\%����'N�~�o�#�D��X��vGz�A=��@�{��%��5_~�� ��v�ڇ8����vKFF.����\��8_'��ݑ�Ӄl﵁�GPX�x��&L�k��S�2���.+`6�y�5 ���Q[�"��!�Sj�*�$�+F(;�G��E�Cf��&��$�<���9|c��e5\� }-�*EךۑsD��A�&n%DM���^Z�V$J�H?<��pR��Y��%�m�q����~���Y��|F�A,��/��R4";��dI`����GY-��՗���.r���P��ԙ:y��4�>t���{�P���h�Nh��Ⱥ�*�4���	NE���o�}t�Ŧ�m�l av����ڿ�w�5,Ͼ���	-k]��d{�GgTr��ᤱY�x-�;�%�[�$IG�Bs.q�����d��1ߢX���zz�t�$��]I��#e��c��)7w���Қ0K'S�]T~l璘�*�� ����XvA	���k\�D?�f����O
��e��7����?%XSF���D��>J����W-�X�|+�&{x���?g��a���/�	%u�t��qi�=���fn�4�w�^m���TxE[�����m/���^�<B�-X���_�b��|W�-�Ӏ��S��α�iE�F����Oz�<Q���c���:Au���Bń]с挪�"e���`w@�oXϙ�����U��[<G1Z���o�}� ��&��p��Q���j���d�_�H���Q<8���L����Mf B�3�u;������\�dk8j��?_�<`*��W�L��Y�r��U�Q���\$��д�ׄ��ּ��mQ���7����1͏���/�� ���e�J?{,0p�V	���'\¯Mg\~�gHN("��JI9��.�~~�<k����3P�g�_[������"tmG]&b���a�?@3Ws�����yN�G��_2�l0�fs. �S���姾::�d'Z�7 ��w��;t�?h7��6 �V�q��+W�Pp[�&�7?E��~���4۳�`I\m��ĖS�-���5p��x��7{^��1����;�Y���*I�{X��� �Ph �:Y����S�dB6�տ?�I�%�x�{ ��`��p�J�/]���i��2�r�|�a"	���q�`6z�7>�DDQ�M��3�Gʐټ�6\�>�(�Ff��������7�	���.���k��S`4��CHZ+�� �:Q��D��h���|����O�رzO�rE�iN�#!L���UJ����B����7��?{*���Jav5N����+�=�w���H���Z/j	8�ý׬�S��������Mp�� ���"=�����ӕBz!i�4_�rNr���K^��2��D��[5���L���:y^�3.,�'�kU[e��\-�<R-󢯻|�_����fB%���d���y}y'�2*-�~�{&���Q�`���7L�m��䋵�%$K��>/͸ 6R�>��a#U�̕�\�\����3	R��y_#��=KLx���E�TJ��R}("�� KiJc�dy6���K�]WBE���&��q�8.S<�iᙽ�S�28�����҅dl_�a����A���{���!�#��)��gZz�]{ir�4�yȁ0�����j��4���A}������̞ǈ'+�L{�P��X��n�-��d�F)髍�#B��̋= ��jM)�����#���Ϊ��O�iĮ����˻�m�k�Ւ���y,�|�Ž�>��PX[3���r�k�u�Z��c�9	�?!�Fx�D�7��g���P ��ݛ�δQ���7���G�'2; �l����r?�S)�Ez�Ǐ4�t~v2���x��#ہ�鉋��^�rj�}5'���g�M��8퀦T.���	�.�Y1�vCTd�̣>̚�X�tfdD���)R����7+{�!��'-�*VnJ�|���y��ǭM<��3���s�o�3%1g)�+9�C.�=�J]p�@Le�H���<b-2�6Q�2�(�F�º�������j<���=5�<� ���k�`�I���9O���Ģνk��r8�$���>������GȱѨ��ʍ����uH�Y��F���ͥ��J�&'�[¡L��µL�
�nw�7Q|�s�C�DČ|C�V�c-tTyXm%� ��X���:�n���ݞ�r-�J;�p	��SX��ȵ�Z����( ��袚
��5K��y<�r���,�}�5�3��
� B塛��X�8H��=뎒U��2�����*��OY��ntY���$�Fj� /x��L��:O�*X����Ԝ���ɫ�h�9-���B��t)Y��1r�i��NO}��ww�s&/�����K$�ϰu'Y�z���N�w�h_߭��6����n̩?$O�Xr�P�k�wq&^c��ﷸSNŧ���!�j�m+s�.U�PW!x�&�G�tFtxP0$N�Y��з4����A
��'u���#�a�iH�����r�ړ�5�N@�r-.�%L��ڥ�*�eX�`2޸�1�ך����[[�ؼ��mT�Qm��x�X �S�սw��~���x��@ٳ��bM`��Z�0����H=z>��Ow~��e����2/4������c��|7C�6��a�c�F0G3��Zt[`��ӧ�-6
(-� �y�I��H̘��3��t���e/2 V�En���Y��48����^���S�'Ó���3�-2/ƌn�]A���a�FŢ*H`,N�'�"��`�:�d� fh��[v�j0~���P`ρ�ovg����ؕ�o= 7u;�&E|�of� �"0@%�u:f�������*d[���KM:�����ysc��T)�l����,V1ch;bU_��w��4a�.�H��; uuE<@�B`W�H<���[�cB)�	X�$3̠�`��v}��=C���c5gH�ᐅ�ߵp>K�,�+ި�i�u8��z4��,j1ن�Y�\��d$8a���T��_1�v��9C�޲�ĵ�B���z*���}Ӥ��@��ѯ��k>���:�<(����t�N�Bc&��?����LAM���W`V>�xy@æ����K#�H�8e��X	p� &��'X����}vR��"z��`�mB���:���:����Ԝ�N�����b�HJ�ݪh��`�c�۔�^Mi7��6h���.Z�g��T>x�������U�~O_ōЃ�A#c	!�#�8�J��0�� 1�N,3D�r�Lɽ4�(P8�n���)3|�m��V0�mK�}�*������̎9ҢSP�d��y�4���*���
?�*����,�����	Mi ᳺ����pS�-�j�zlj�c�Q�E�Q�.�|C��޴ý��טt�=������u��L�DZ�\�0��m��ֻ��j}�^ͨn�8�'[|����$6i�7�*]��VhÏ4%E��/V�a6�e�����>\0�7��3j����1���]_s�Q���]��c=�2T~k��g)�Cd��a�D��$e���^���G��*LU?S�	6`1�.�/�����0*�ۅ�SpF��-�1 �e11�y�.=Y�Z�V�&:E XR�8�������Z��%���� o�0!�H�SR}b��C��*�ֺ��=j�)ǫ���2� �
/��T����W:_�J����X���^�reV|����&c�����ǃ�1,- wB�[�qw<y$dI�e'8*/O�(��̸�-2�tt�GEcV)�4�z\��:�`����s&Hd�{
�G�U\_<�7��㷱j��A�V�J�Z%3z�RT�p
As��FLms�����SU	m��/�+>z��F��a\��s�H*)=Σ\��}�偊q����_�;��!q�?}�hu��_d��k��G� ��ލ��x����y�|	�\!6�z��kJ�K���p�\؛q"\�JJf�q�q��)�A�EӅ+*���N�ᯈTh�����v_�$�M�ցM-�<Y�]�����sn�.<�ϔs�8��ZY�����+�^D�����(+톋_f�iQv��w��LtqE.a��PhZ�4�_���^rf
y�Y����t�|�e�uU������\�yg������>��*�;v�>��*`0�:I3��k�vX?��.��ȉE�yJ.�Y�q0�����5n�"s!,o�gӁ{�3�I�H���@آM��+��:�:�H
�D	Z��ystk�!6�2J�������x��@�I�}��d@�;Jdid�5}Ҁ;#6�arn�7�3S%~��{Fu�������6<A2�06�O���UgH�+:���[ڬ��Ϸ��N#����5j���>xj�$�?E$�<nyCe�_/'FJ'k*U��a|x�x��77r��O�A��Pk��_em�$�mhX����\\=���G��~�jm&[wϖ*�7V������E���g��s���k�� ����
:�B�zRSz��$��)��Yl��VK��,����һx��#��-����)���=`�%sH��7?��5�e�n�BrT`�,�߶)�x��]$�y���)�������"Me�rG�s��sY	0��Ϩo����F{��t;�d�j@�ڳ�n�~樒}C�lvm=�e�E�?��tO4�*z�|��аȚ�OG����DwÑw�XoA��Rd�Mg�bDc��t?2j^���8W�������Y~l/�4�4�@k����w`�RK&����4RN�P��T>����rw���K���CA�Zn�eq���׹c���|Lz����' �m"hg��8��WO�J�������|�b�� �P�
�6�q/]�=/SB�Cv;eE�c�bJs9ו[Sj	�����k�$��)�b�-d��<���:�-��ӰWg���B0�(���sF7Fozb0��B��Q��GX��p�X5�jU�Oo��$�����E��j����&���jcP�Z5�b���`1��EA�Y�=��R���׻#��K��KL� jP�Н�cd�����1kC~�ܟ�����Z��E��O"��Õ0��7)z+�-67s�vR;��j�j������M�zP��{�2y}���i��&U��
�<]���G�'�֖���
t���|�$��p�)��j!�&:�c��X5��t���﬷D>܃Pw�DL�vҐ���Xk��A q#�<���e�l;�4��$E~���wk�Hc��j5���,�n��-�Ěm����z�
�>c�n��^��hjOТ=��Xf�2jca���$�&�)���\�)I�@�:��� <B8B*�8�+z,��:R�2z>��|���T����\{?*L�HKnF���HKiIh�f�IÇ�4�Q/��,O|嘓���[h|eI�;�I�/��g��h�Q��^�S�����I��t�Ct�:�v���1��3�t7i䉇� ^�� fa[=�l� �LSnw�T��8@��
�����}ƽ�Ȋ� �>=Օ.۰��=A���^O/�#�i�����&z
P\���Tߕ�޴�����b0�<22s8��v�	s?��H7�ŖM���J�Z]Y��dM0	��%F�٠sח�3W;T��GU u9��w��^��yqkse��Y�8�K#��u��4r��,��\a"V=$����+k
ٵ�>Wu��t��jDM=�"���Gȳ�i������tk�[���c��*�B�l���!���OD�-��Tp%uz�����q
 z���TĞ�H�r0H�J7�����q����	��a�sUw��E��04tK����^������8���-����~f����Tϫ>���^e�率nL�Ћ�u�:d��-�.�?)|w�k��e�m�b�s�"HW 9�V�=	e�``B��[bs��Lx��mE>K�	��C}��r�W�Y ���x@Wև��<*�f/�liJ$ � ��8���I7���_J9l_gW�{�L,�FY�s��<,:�N�1H��m��[�& ^;]���0�����;�&c�A.e��.�e}�
����۠M��dΏ��1�q��GČڻr.�D{����x;���ҩ�8df+�q�jTUȓ&/�)+�q���ͅ�'-5y�(r'y��%z�I b�}w���ȑɗ�]CЂg�~
����~�d�@����5N�扽��@�� ��#F^�f����:(�?�+Gj�YJhd=ֵ�i�)��p�AH,���ܡ����
f�B��W}�_�Ax�ǒ�F$J}�ҭ�����;1(�[��v�k�sz�^&C�n�Z�*������m�:�t�N��C��������G�T�D�Ɠ\ZA���hw��f�t�)jV�2׼��S��&��_��M�0k��]��U��@g��&�*6�������ڧT��݂�iJ�c�ǂ��4�9�dp�\��'Q��2/	����%�G��jT�j����8���pZw�-ˋ;���,]x�D'`=p���+���c�ZSP��W��*�׮�?L`/I��gPˁ���+�#�P��&Q�6��Q���mI'���U����yҍ,2��G�2�ʼc�'_�2zhz�\���\�@��V��z]���SEt4���QwWt��*�=�18���7�-���t��YDufU���"������a�O��݀��mh=�|;�|�ђ8��g��	��%�̠v�I���n�q���9)�#��r��������Iu��+U�.����E[@
��`��Tↁ^RA'"��8��H�;�N�?L2�{�~��PW ҃w��	LVIjZ�����f��n�������wX��jk���+A9�v�S��5����3GAfE�[�~�B���)�r;�Ϣ[��)���6�8	��1��<9�ƵDH�M
=v�3ܡ�]�2���(����`L'�ݦW�5�NT���R��P<a���e���J5.ADJV 5S҇+�[��0!��p������6���U*��Wo�^
a��o2���)�OT���[�Nd��A��pZm���J|4X�˸hV$���pk��`9�,l\8E;��9�'�Tw�R���'��y��`W��˄Y������Nw�D�Nx�*�f�綗��_���ա�
��/5����&ic�k��^fk��P�P��q=b}�=��YY5��Q�c�|�s���Oy)��Esϡ��ޅx�Nrژ)2��T�qsNwG���ڬ����q;Q�*Șd�#{R\e��|�U���e=�_(d��`o��&�x���f�t�����ƣ 1�ܻʕC��� IF�	EDڷ�gO�Cd�����1�Ѽ���'��bA�[	<�1t��pVO�rb��u�d��S�Yb/m�L�qp?�C�R�a;�����K�o
{��\
�kN3�_U�����R	�9�2�e�����;���������
��Zc�-G��L8sq�"��pfT�Aa"���� q����)� �,��Y|���n�t������^���3��}�y����@�<�6����4���Cn�ź�/Ab+͚�pynk�m��c�l���*/�)|�������v��=�4����׫�>��X�4��}u�w#n�������v��4���]��z3�z� ,{�Nkn��	k�1�������2���mE��M���x�b �s�a�R�wIM����ҕ���P\�J������~X�R�X���)����jO�3�ܒ������:aъH�h��s�}ҿ���k"H �N���+�Q�o>^-N苅�*<�V31��>��
��cv�͋�H&����0s���3P0vC�9� G�6�T�\���΄A��%4]�N"��d�ء�(�<従F.����#��_6E"��n��:$QW�.Dt�����_�>NB�av���3�6�|�� �1�i�[��w�%���D��u��B�AGu��5�ñM��»|�JT�,�޼G��s�(9�4�@!��{!����ɇ���8h�(��^�޶��3]�>���M�C�D�x�|Ψʹ�>���*�:m�~�� B��^�6 �}�������)��E_�$�9����Q�������k(��k��y���L:����INv�b�¸M��E��-�Q��z7��BZ�P.��rkژB�������`����#󟣭k�֪Nӛ$o��g�0y"@�#g�l�:V+�;�کT6�}ˋ�:7�U9��@[@h�tp�����;��#G�Rg��r�q��ψ�~u�[�I�_��]x��x��k���r���G�c�.�j)P���4,u VFs�V��>�zՍ1����A���㬕Q-] E��7C�{�M���&e���\&�MAA>ôv�%��������X�F��؆Sr�9u�/p=�ml�S?�z��u�8�D<�̾J�*�5��X�~+��N�ءؑ����=K)�>}��^[�|��
��`��a&{�Cּ�P���f�����>?>�9�W{�v�R�ZyNSȆ�/��,����W˪��	>ٺ��Ń)_�S�L�qX�0@��ރ�J+B�S�jw�%�����h���D<1�sg5:��m�6�7��N��rC8&�;@+�ʑ��
�8x�%�)���y���Z�$�k/F�hR�H7�
P�ۦ�_zN�3(�<�M:�k�&P�_Y��n��P�S`mmW�ğ居6Sj��kRӧ���Q	��#op��0z���T�i�Q,���c����V\���*3H�Ĭ�WBpk(�:�6���!�Pz|G�m�y�)�v���-�>�=/���*W@a-��ק�V-�j�Gw�yI��(���8�Չ�
M�0��E��@�<�r���'�����N���8\�[�b9�t�fK����⦗B���̋�rPbH�j>M�)���4��kBK\�w�Eۑ3�pv�������u���h����5*��"1��:�!����Z���m}L���ɢm�1�
��#���=��P�dtϿ��	�2�!��~�ˍ&����z.ޑp�?�# �xv�>��
}��#vuh��j�&���w�3e�.�h.��8�l��F�=�Jғȡ��4B�A�-�ky#�_�_ _,��0!5џ����\�d�k�}�Osk���S�_�� f��e��wȌٗ��sK��Ē⦧/��������3e��1lu7�:wU����̦�V&�<�1jc�3L������+�n���d�|B��}V��Yta,!�{}%'ށ�*h��WP��W���F�d��Ò
�_׿�"�C�мȦ�G�����u�a�@p�;?>E�ş}�^<m��(��Ր=�u�Q����T��i��&%�b#\]qmm�r�A��>|���J�:JG�t�'���Ē�3&���_�o�D�A�hV�M�ys��e�E7��&���Ѿq�ԫ^��.�SF�T7epYcq��U�%J�X�JH�_��jɍ|6���8�~�3p�빎N ���ݓ�]�F6��ȌD���hR� ���j��ߟ�oHj\"�,4��`�Ga�L���qҢ%�||�˅Dڇ�+�QIY��q�VD�$;x�o��@�C�c�?=K� ?�M�Q�ں�5�	S���+MB�~"�N`���G�oM�Za=Rtc���Yā!���K�b�A���9�ű�Aa�o2�-����@t9K"�h���ަ��U?X��e�v���>�ΡS�<׭���a�5L P�z��U!%Z��&Q%��q���|�	gJsI��5y5|�Z�u�+B���q2�g�P�t?��_1��@�4��-`����֧� ���?��&'}��~�8���&�N ~ 5��;�|�^De��W������P��~�o���D�k�Q�t�;<w�ĀЯ���2.�j(�H*���k,���1��g}����Z����-/�K)�����PD��k���!_p��_���|?���m�C.����`L���*�Z���
�Z"R�L3S"�٫�]t7��>�B�;�����K@��,�Ōw ����=X
�e���m�I��<࿔.���h@Kӵ�Ofl���l/.f����M�@��_�ey�xqE~��{����h�O�u�;� 
��ڪ�!'��A
�캣��ce���I�rT����x\㤋ݔn�l�0���]�i4�R;~f���t=�jQY�������&�	�|y�%� $� ��n݅-�[Pʆ3Z���1�0C��d��r�f��W:�)z8�P�Z[,�Qr
s��C&�+�i�<���ө�,�AN��s���Lɡ������rp/���� δ �BG�-��~��y0Ɋi	i��6�wI1}���;&͓�^�L���7��/O�z�2��.��4kpOe���������Wג��~��t��p��OL%�,֑�D�ء�׳-9�7Ӫ�țs�����쏿5#���v�Z�	�ى�	�X�[��_�����V�ސKP��g�-^P�V �������$��aٚ�2P��P]�W���]�S��N�Y@o�{60��h(�xKX�ŗ����t�g�2.��Ŭ���M�)�P�h�|��CHD����]�֒@Aw�`��$�J.��vג.-	�漌��$I��u\���i��&z��f���T����0Vs^ _��]Z���9�C���W��@-AsJ5��V�G�̾�mZ6�&0O��*jjO1uC�ۥ	:�����B}�N����v�����R���1��$�T�(�Xn[i�Ϥ�@2����=q�(*�� ^v�I���x�;h�v��y3�1�vK4G�VR�ͪ��"�f�ys������W�1 C$A�<e�Ń��^F��g��*R:�2�� '�����l�[b�C3��:�f�'y�Va�m)Ʈ-TK�͖էH�vF=� K@�tt��f�+��|(38�Cyw4�9F"��Q7�AA4���7�]d���28Y��I����9F���j;�m�M�|~g��%�` ��7_�2a8zW���U��w^��Gc;&�4L�� :�����े?w�W:�"�>��J�8�3�ȚSS��3�hd��:Z}��e��ҧ�pg�×e/������*Γ@�|�>@��;��g�cr|�(��ٖ��Ǯ�""X�����e���9���~r�'S��Fc�PċiF��.񽎠Y.�8g��K�\�F�9C�,�v��)_�����o-�6��|���kDv=r��ހxiR:YxK�/�7z��l��ʛDm˭v��Ul�^��>��4	m}�Ѓ&��'8��K��̛��0�����/w�8G�<f�a��f�����Z(�זn>���a.���0���]O	l���g�o�,��Ms�w�������|�/�){�/����Q�{N�q 8��q:���R*hQ7��Q��J��s�������/G���T�~��6��e��)z��Oa�Z�~�e�����y+�u텻��Q$��D��Ճ�G��J��7��ɭB\1vq+[`�ς��V-��*ɢ^����m���p<�No|D"a�q���< �`k�NqV���ۨ���e�����"�����I�؎�}C$Z܂�%�mݦ�pҟmG�6���\�����Mlv��K�2#<gY��?'`�����mCM��e���3�YSg�eL�E�W��)wG\��W9%�5�Ӈڛ\��;w��\S`@x��� ��tE��з�>���fR���B�w���Fd�I���KL&*�ӈf1��G�!�+���\hb���B�-~�̱C��'�A�A`�"���p`}�tN�F�C�>5J*��k�O�%�/�É��4N��C��eZRɠ�U:⍃���8���hԌ�6$р�}�h�6�᫮���������%3���H]	ťg"�� M
�.�^}D�M�i0�M�=�ȡ}L�)�I9�𖏐�y�����q����!g'�����X:�g��6�j�\����"b��׶fm�2�A�mB�2�o�q+M��2PK�T
Ne�*�r�õ��.���.���xt�I�2*���f"�Ғ�VS H@�'���%�V���{�JZ��NG;D:�w��Ix�ljD�[߮i(t!���,;�מ��:qO����d@����z�O�܈��� ]�o��U �fS������XZjPX�l�qi�}E@1�c"�,��Y/�s��X��6�O�r�ը��̽x���w�Yz頚�i+Z�s��LH���y9�6˽Ux��:1*j�m�uP�w��_���ad&p�
��>G_^��ͼ=V��ow���4y@ܿ������z4Bj�o�A]���1n=�L���><%���&}�xX�h�� �7��	;���B��A�$7����އ�ˡ 2.}�;�"��Q�ͣ�/{��`;��`4Ǡ�p ��2�^s�v�S��^wY�`��α9A��e�wR:�Η��nʘJ��"<r�⏵5�ч��NWJ:����G�$j[���ұx%kq��c�
:�O��V��A��lܶB�e��L��`8-6�P/�:���U:�tFxt���h[K�L@�ӹEXljA?˺5a5��\�����4*��P�Cqh�p��q��p�����ٛ�4���*�]����`$�<�Я�\ޤ�`n@HH�|��Tӌ��2ַŞ��?К��[�t��<f2�o�3�9��� ���jM�Mq��Ih<��+z" �m`��f�B�����Z�!iX���_�WY�?�`K��9�P���I�,z�g����6�(�;�"�}��c|�:g���h㫉�e��H��$cyo):������轃�����u�2����F3��i��+�}�b1��H�7z"V��ܗG�������ix]|f���I}|��<����m�r�a/"qaKKn�9ߛ�7*��	N�V�c�6ķ������������\}�i�B��K���}I]�����%*�^K�Q����D�?w�Q���=��|��	���;ѩ�Իo���MW�z��h�=.5�|�^fʐ/��/+u�m�*����r��=�·�I+��m��B�ѣ<���&�֥#������%j!���E�W�@t�|hZ�a���n��1|�eUuTqj�RJ�
��E�D)&�1FypZ����E��(T/�eV���r̕�Q�l�([�(�:�W�'vu������xm���
�����X��痒�xjDq�:k�� nX$]�F�|�/�Cm�Ĉ�r㪶�3ɏI|$�0���1O�^N�G���}��ic�-J���\\�§+v���jȢم�]�5Xa��PIb�n���wkz+%(�e�j�� b�}f8ݵ�>NR���>�m�ek�P��m��I�${�џB���ę%��ต��!B	��~u�>��	k�=b#?��!�bգ�eflA���I���Ҙ�|+fAc{�dM��DM��A5��x�n�|E_��;�X��oD�6c9�곸p)_�S�!4�n�H�"�,\� YН�ܦ:T��mEЕ\6Z��O3��k����j@��t��6�]�Um�oŧ��7�>x��43�s�u)Xu��F�E��fs�\�/Lھ[��=}���Լ��J��FH�>� �<,�XJ�ڒR�ț������R��Q4k��F�-�����:�t"��ѐ6]�?���/�߷�ҭ���."���!��:x�j�����I� 4���tI(ȯd�[0E���01�
�{|2�+
�+�%��A�\i�B-��?�,"�`�p�[EdL]����e�4����#�m�Ņ������I��т����o(�Ԫ6N�ِ3W���J�!��rwN���&�^�R�ϩ�F�i�4њ� '�yX�c��N`����1�i�U%%糩��]�Ք��DA0	p��G"F�����9۞4
��Cw?��gρ�oY�?e++]�?��"����K����4:�X��)n��B,݉ɣ�	1����;�|���	V�V3�\�2���B�����k��f�XZ�ʖ4�266�gq��ç���� $��H5�:
a�����j 'Nυ(vJ�E�l�Eޤ/��� ����}��֝��Ln�$�v5�cL|�I��Ú���l"Ӿ,~`��l���`C�j$"x����n�~�=�l�@��?$�ίA�9,|F�1wBZk�L�� qF��\3�{U{s����(����>�yW=b*;.����v:3$�GI�����X��(�|xOzu�u8f3��X�ר�S��dC��0u��JE]7�}� �ZݑM~uT8��	e����r�#�+[�TFŮ��'4x|k��O�:�f{g��$Ø�6Ѓ��DL���~�2ʄ���q�E2�Y.Z�X�8�qs�_���3�*�t-F��M �w��F��+�%���
�2\�����ݿt������I)�D�K�gV�{\>s�=��Wf�9z��+�7���b��y7����S�h3K�L��rh+�(%G>e����D��Ϟ�c���>��Q�*�l�,M�1��F0�ӫ��3R�ҿTm�s>��ʭ{�!�%Ԃ�.L`"�Y��
(#�='�`�+���Z�\�y�U���C���,_�˶*�F�n���("�n~Ӎ�8�rX�6H���a.�lm;�c�/�xYJ��p5�H}9����A�f
��T�C��.8������S'�Ũ�s���ڸ_�s�"	��-���̜�Q��|��^+�Ϯo�?�޸��Yg�c�EB`�;y��J�������Sm�X=n��[�r���4$������m��U؟9'j���9�2�f$=a�۽�*����:k<�aI�\���?֧�ıy�����]�b���-��bt�h�+���Ł�w[4�țɰS��m��wֿX�$�h�������\Nu��]:�y�~��b;4��y��k#��81r�&��)��Et=������Ӿ^��Y}�,�c�;����o �xb3��n,�R<���/�􊤹e,�Κ5<�
�ǏcxJ�xK�*,_��f�`B��m��,uYw���?��#~.�7	5��{��eg�����r�D:v�@ܢc���M4��n.�5۞��8'H�{S��s+�up'��A���cc�h�:A�������h��j��2<;Um��ώK9��h 6��4���;1���ZC�
�V<�"����z�g�R@�~IW�?�y��*���� � �����	'�@&Pu7.b����*���P�Oy�n�U}|(����6��AR�6�_��;�%�|A,jNwO��5�rG�'*Rk��ƽT[f���5)BΨ���H.�����>���EPQZ�g'`�p�i���z��%�~T�Y�����aq�ׄOB�}�5	0!�1t̙7�zG�~�
/�EUD�_�~�ҫ �j�c��(JX�
�U����q)��F�W���Rg�k�v��gQ���KS�S��g�bj�� �NI��]:u��]������cE���}�
��>�49�B�7�A{Ė�q��z�f�ݠ~��2�~;�?Sv��
B�|W�wr�r����:���
�Uv<`g
�:�ďkpp��<������r D��
��:�(��P�"$���9d����ݕm�i|�MՏ引�j��zhय��1s�X�2��i��o����R���,�7�rY�T�<��d)��wz޸l�'g������sO�����y�E��n���AR	��dN)1f���BS����j:1[�����5I���b�~d���,���&>#�=2�t�D\��h5������$�D7�>��Y�ϖ����j�L���j$�!�~������:�L���������Š��������	�a���R�B��X-�=>���Bq��i�W�򴭹\cU���<�s֯�<�&ԯ'H&�m#����Q3zD��Fh�B�ޝJ���Fu�j}@S3V���u��CD��i@c$-����y*;A�t�::!���]�N�,��eQS�3OvL۵����43t|+`ѿ2+m����)�z�\Ft0/q[����G�l2�%Cxmޯ.B���9�,��"��C���ֹX�{�H�����q�-��
(Y��x�/�z�o9a�A)Wgd�?�5�EJk.�_8^O��!a&�إ��Q�k5�p2��^G���Cє؇��h�D"Z�٥�K؇�����Z�Ry�88TB`d<~쿄?��kw�̟wwn������K��U�+�J������e�F�'�3�֨�g|�C!G�'m ��kG�R2[��!�c2��	�*��"��9����"��W�U^�`���G����a9��.^j>f}-�y���d�}=3�'/�si.D�Źgu�V���N4���㇀�&*oC��MǗD`� ���X�n���3R�z�Ɩ�Z^u���������k�� !Y��c���m3�N�xg�2�fU�z��Ó�v�Q��۪��2rv�8=�V�c3�Ĩ�(�����;(C��#r��`*=f2���Z<u�Ņ?=�(Oڌa��q��X!JD:t�H�ؑ�kj��fQDP5 jr\��k�Ú⽾	�nyڅ��-�-��㿕��bʼ6PM#�q���6:g�{��dֲ�>J[��sћ�]-�^%����5C�=ʸ��N� AWF����|֯k��c7��X�pD]_���5~NǦn���ᰊ�EV�4��k����D����c�\O����S&��R��U�씡F2EV�W��m�pc�^'g�^�OƟ7
e��6u`ϴ��*���<t~��YK���l� ^8��J���W�a�N����k�l'�>;��n���^���dvVI����-&�#u���XD�2)�� �f�31���xP �Ҿm�Tz"�\�0s�����w� �T1yǵ��v�k����K�N�(��ɽ_�w�(�!�̌���A�d^p[/�x3��eke:�3Yb��Ks�����I�����
2(�D���!]~!�#:�
c������b�0ۼ(H;� ���h������*Жc}F�Z E@U��F�1H
"N@O���/�:�z�o�S�k���zR���l��;�mf�:=*Rx�nۃP=/x���S����6[v��I:��7T[�~XY��K����4j�,li��!��5�ٟ�\��a�폵����y*z���D����<ͯ����&���w�jH\xxZ�Olą��"�U����Ƀ2d�vB�j���߱-W<	���ᐵ�'�L-GR��
�F��ɇ��"LC��\�ͯ�U�nv����D�����ѳ��е�sR��[�Q��@�n��"���X������6��F�ا.�R�Y��b��:�\w��yw���������I�b+�1*O�� �gG[�����������4u� ��E�!P��3�ˀ�����E;���z?o���³`�<���=�&���z��[�O��~���uhgG;ӄJH���X���^�ۉ�$�� �<�2?w�J���Io�E��܍�gx��(♲k
x"���ċ(������1	=���7:~�^<**��r�]cy3E9����W�aO��A�'��}�?�����d��r[?�^�,���uw�j	�W�����LR�N�b�_�ɱ)��b�	uo���-:NR�^��f�����h�rK�i�$¶bw�v�4N�z���_^y=k����1z)�(�7��	mì��ƌ���w4�����H�y#��@*��
���Oy���)#}Y'׍��[�d�(���4L�v(��ν������nަ�N	�]�Η�K�ւo�7ֹ����'���1%{o>�Qt>���ǟ�@feM��D���v�k�H1K���#�Ɇ8� ��H�$|��Ӹ�V�b��tA��`S(�hYK`W.�'&��c�����+���K-c�E��F��Ż�aŌ=w>�t�rAۖ[AXD6,�f+e������{C�rM��l�Y�w�����w·�J��`�D^2�&9�]XL�tX�8z7n�?�@��6K'뀫t�����tqS��b|Y? ���/��;�<��9��͎���W��Y����x�ru���:F1���\	���{H��%oJ�gm�U>�Tv���g燶'M`�oF�yt~�Y%kWI�����,�����2Vt�_�� 7���P��3��`]�rԪ�X��2���TjI�\f!��MP�RŮ}����g����W���\u�$�W�g��8ޓ ��j�C�a���qMo��Z"���3�v�w�o4>4���� F���V=x����)w�xE̿�7#f!���"+�jI'V��}Olm�%d�W�Ջn���r�~����#\�8:�kE��}��8�Rc���KDGtj6J@��;䈗5�S�AKN|ja�|,���t��{�;����/vԝ(�@3F���^�b�wYa���62��Y$����A�,��!C/��< iI5��Iߜa84��K�m����m��<�C��w��3z� ���G4�D�m�� U&��й�m'��J��xc�<��OL�\ѿ��S��;�+e�'�W���yô�������A6AD��~Մ�G�&1ʏ��Y�k���c�Ny鶔_�5���F;��������HO5�_����'ӏ��
�+5�ɑ���
p�0��TST�q��4�ς|BOs�q��.rg�t�S���A� i�r�N�Bo �;����R9���<���U����v��Oh�[�j~9�<2f8dO�F������䭘y�(��*X��������2��Ek}ː�1U��&R�,�0�M��]�1y�0P�⋑�I�wO>��1���Y�;��vP>o �K<چsJ�@��o�6�Gǧ�`z��򘮅X�F�|���̽KŴ��1��S&������Ĝ��Ĥ�*�1m4��\[
վ�EG��_�0$�0���"���\QH��c��`.��ë�TR�7*A5��:Z�*�_���Id��j:�_L9��vGtUn�iT��w�l�lO��3���i�2Gf�_A�=���!KJ����m��Iٰ�����-`����$�3C]�6�#?�4�H��"fpAX�	�(��Q���^���D��D�ގ{��`�Qf[�H{D��W��zG�c�j.��bh"��C|C�=�w?��:A^���˹�>�;Z��
��Nˢ��'�����_"s�{f����J`%�y�|����'c��eb�6��Qf�#�h������h]t:�bχ@
V�{n/���ޙd!�K�<9_�;�D�o�LA���{�����{�=Te��o��_��B�D"@�l��O��y놇��j���
�����x��R�=__�~v�[OZ��ESb&  ��y l٠-�'�/.'�Y	�bꞾ�_THk񋳦�/yO���g��C[��}���Lϱ�մ�pJ��<XE�dK���@��x�HNg&Q'`~6Ɗ�sމtlZ�*��;��&��O�d3���$�Ov˶��NҌ持u��
WBy4a�z��[�����������Q^_��6���U`	�0��6����N�D|��!�� �&�Ŧ��$N����S=q�n�����[2y�f�M�}M�5$gOX�D
�I��X�D!	�C	*R}^�H�d=V��WJ"�;t����Ԯ�����T#���Q3�|�����ߊ<��/8�>J�������#��8�eR�H2�_ֳO�v�d�mc!���Ѳ`�����WG$L	ڒZ��W� )7�8u<���'�-�w�I6~	��>�oI�=$��76�����dQZR�:ȍ'�9���p]A��'a��+��i�Y�����%�K���uH�K�-��9�8�3SP��I`nJ���bD���ʨ�l8��6���uI0�2�)�Y�ڸ����h̜���F�E����J���"����/�UʲF~}c(���m��Y|��P]��*ε�$*W�-�V^n�~cS�������+K>��O���4�N�2�����L����F����i!+6��1�d�q��!�_�մm��_r9�����O\��\`������u�R�3������0UR��*�����C#�"�l(����}M(�z<3�	�����ɉ��i�| �n�1�:l��_�^���Bń�̠Tp�#ӁLg����$��i~�	�;�)��������:^��!%5v�^��&#F�|zj?���G�t~��$�����/B�O�
}��/b����R���51�`oj֓�aO�=���K�od��Z"z�M��o�}_�1o�^q.n܋M�#T�3�*1��
P�9,�xI��@�eBCxe�ݵ�p�5O����\��	�F�p��m���K��f��Uܘ��D��N�54ա�UTKR�kž��T�l4��#x���4E�);���+�<?�6!n5$�GT�H��Qi�6�<�õ^L�x����@\;d��� Ȼe>��Sbc;x��me'G�E$]�3k~�y/YA�*�-�W�Jo>�nA�D㝍�d�~��%��*L�ڡ�c�����%�8XvN��K�$�$�Zw
�F�[.>�Lb�����1]����ޜ1Σ��|��Tm�/��H� �ė�:#HsKeQ���N��1�q�����_���s�+�m~�H- \�!�Nu2ge�~�_U&���	�"����#�M�	<H�{�A!�X۽�of��c5`�Ha�iL�g��0�JYDq��tµ��7����hwk�~�{��CG�83�<���q��K����;=2+/�C�\�a+"��e4<����3.n�	��)������@v���~��.��0b�Le��S}���Kg?-=��I�^}�L�z��WF(��#�	j�7���2� �xv�1I�"G~,d��BΤςZ���D�Q�����Dk��ݍ֢��I�M�.bYu�R��mJޏ����ՙN�8:�V�)�$��ɀ�8צ'� ����`�ju_Ш@��y�,˃���P�4@r2�m�b����Su��`�{�)-m����`��,�9W	��	�ݺzF�PJ�<�����N �M�p�b�����u�M%gs�my߇5{�uZ"���da�Rz��VF(h.�����{��Ͽ�	�~�g��>6!�fB�-�+�j�O�+��;R{P�Q��93�◹���?�����qe0T��Ց��+$�f�?��Ag�',O����*9��ou��t��4�Ԁ�D����;���dU �z��7�2��cԮ���4s=�H�t��`�遐��V|YW� ��6��uI�%r�z�jp��a�����7�
{C�oN�C�����k��"�-"���	[�*M/x�����o�z|{b���o�����.��G7���x㕛�\���t-�oj4s��&�ހ%3�jE%"��1Ƌ����)=X8*bΪ������ӌ9:C7�z�����H���Oء�J-�3�Q|��YD�P�����榡��~�p��]K*h[c�!�!�'�@ӵ�y������D�c�+�:C4޴�V�L�6�8��/[(�r�#�����N��u*���AY"BAN�e�إ<�/�2	���<Y������9�T��i$�(!���%�%��_���)��ȱ���'Vu���ud"�Bu��Z�ˊ4��ׁc�ʂR>Õ0=o� 5�:��,����%z�i'�.ڱ�x���r;XSs�$̓^�cd>��F/�+̵{�A�ӏr^,װ�悞Q��4cg�p���6���+��~l|��Ց
p4��� 5hL���M\���/1���x�eE�o]���W �p|�Y���JA���_<����cj�Z�]|NHq�!V��u�.&�U���X�z&�R��7,�9Ԧ�x���m�qi/����0"w!�p����#�r�&�J�>؎4�dEVQz��r�#}���6�½b�%����
�ˍ�]xi��7���V���+�0�*����J��7�� qY������]�:��� ��~[���q��ܘ�����'H����M���$w��'�wb]N�:��)��5���>�H
cO�J	��ʓX_�u��`�N0��@�C�g�s�����ǢaAI��&IJ��*��@ؗl^t����ys�>fV�>������N�7Ht���X��,
�=�j3�g���ͧ�9��*�������r+_B_'#��t�*��&cs���Έ>}��-7JZ���+^�$W{�I����=�&e>$��&h���@;b=E���]_mB�(B���j�0��z���F%�&4
k���3��N`�,�Q�������6��f����oC�������Z�Y}c���"�-Ո�����Jd3d�=+���\'��T���W�;ȟ����,~Ѐ':(|����N��Qf�9���y��n���K/O/H���6(�K�udnA��1�
9M;OQ�c�f.1w!������������L���H�g�A"�|�c�9Q�z�i�� �߆Ix�X��g�i<a�]r`L��6�܌�#�
�$k��?I���ur)G=��\�l��bE�"X̯C)����5R"�		t�5�G���V���������xg�V��T���Ԑ��t���p��?щ�@���q���g��΢$T�{z�P6�ߐ���e�K(� ZxEKzFqD���,�5��u�aF^��M�;�g-m��������W�_�քB(~QAL1=�v��j�� C���sW��=�/�l��A^A�t����1<k�����_o'Q�an��`6j��E�%+k��.�P�~3����	�)�8�p�D>&ֱ��O�̺l�0���g���w��L��Sw����&T�'��0���9�������EU�!>2��أ�-.���^��ռ�ba��e�};�}"{�|�](7�TA�e4E%"O�-�7w�o#�XM��mތw/kʃr���i.� o��B�mG��p��+�l��{�)Q�a�ϼ"]����u<B�ʗ_s�fU%s�/���0��~`ڬ�nW+m�U+'��Ku�P��:x7T;[ !iF i\Li�``�P�)d��I���$3ƣ(v���w�}Ȑ��Ļ�����e�:�r 3{k�%��"�T���F�8 ����o��l,�hH��g�6�YT,�.׌Z�@l�ϯ���|�"v�z!�넱iq=���]Kh5{���Op�\�2(�N��Z��\k�%�p�O:��xςʠ���� s����^�|��p_�?UR�g����+�����_�)�W��7�ڇ� �ƽ3����۳}����f:r����7�P�9M.�j��'�[� ��8)�ެ`���
����v���S�4�V�����,3D�S�v�x�S���C����l��c�!<�q�<-�0�������`�g�l�-�m&6R��W��-^�$���~	��HV�J��6_��ɺ���`�sP�>_:�]z;5�s6��0J��ˆ[�,���1�z�i�S�����iأ+?\g3�fȤ���)8�����*��QiG�=�+����4�n�;GD�ZJx@/��`K,���2�Z�~/�,�"���HhqJ��z����El�ot�ejꘚ��5ÿ��x{|����Nc!��a�������)���/U��[���o����'���gqo��ZA%sW'
j̹�?o�R�f� ��1��-������.���U��^H�c���}Ur�NN6��J��o�奀K�x��V�ԧ@��G��h��_�5x�	�7ˋ`-͚-������;�Y��n��f(�3EXo��>��i 2����vOfu��7��KE`�X��<��]�;j����rn��k�v����d6=f~D��L��p������T\n�h��T|@�i9& c�첉��:_���a�a:���u�o���x~�g��,���^.�\��V�,��$^v$�D��%���;oJ34��,����x��Ҹy� �r��g�̥����9����R��x��l�����@=�������Hp߰B)�]4�X�m��T��L�'opd�|����W�|����ـF���.�c-R�O�,��+�V+2�Cj�h��5 �[.��H`�i �iD$F!Q�U��E��$̓K�W�g�WSCu#[�?Z]Y���w�!Cx�>O����hw���KQqn�X�fR-�n2�r��Q�]���օQpxR�F����`�a�BG�"��!���e7�(-B52Z|�����y�,�NQ1c>�v���J�l6F���l5T�CBJW ��8i^9��MO��B�P��P5��X��cU����]T��r�o^E;�nǌҧ
�����;���>���dX��� b�h�щ' @&�W�e@7�I#
%��)l�B�1b�;,����y�&�1Ӈh{P3��|B�-5��3Z�;T�������w��,0��uzo�4g+ke�'�$���(�&(����.6Y��ĥL9Xf�t�fy?Mi���.���ä�R�)IEws���4Ii6FI��M���5�����?�հ�U�Ҹ���4�+^��z��E�����_c&������xNJ�&�1b���g���HN���n2��
�+θ�r�5��`V\D?���`�<�GRz#W��D՜8�@��zC�@�<�0B��Y�^>��q�*�����Z�͛��Wb�wO�}T�4k��A`Y��?�6&�r朒�����1��H�����b�����/��uw�4����#�L���~�4�4/��
a�Ș6k[
��Q��ť|d�'��� J��k��� ����b�;G6���M���|����q�������u�<E/����E������v�9=ߦb�]���F4"6�m�WL$0��7�ꊺq�>���O?2��r'l]�Tl�o���F�U)�[��q�Cյ��C��v�b��=�a�kM<��2���y$�}ç1�����&@�ۭ�e��I��ذq �9e5*
��j�����䅽D��=]��x)�K
9X�� 8r�&�F:	�A��3�<��$�\ba\U�۱I	��Nj��X�P��Ɗ�ឺ��3�d��Ŝj%�H���s}M�N/Æ8�1�y1V�&��ٸnW��忔��5�@�.%\c����簵�k���zpJ�<'`���J�Hџ�m�jO��х2U'e�<���އw�o&��<�b��K�z�q�O��ybg���rYkJ�>I� �:.��C���1"(��+r��،$��$|�C�y-��X����5�f͋�7�F+'��e���Id<��c���8U���A��|^��?�����M����W�Ze~�2�d�q� ���O��-��B��,��������ƳcR.^tr�n66�Y�y�0$ގKhy@D��������F(��@ԑJ�o1�L���"�f!����b|�/oF�%n�A�t77�G5��%�
h�����=t�g���Rx�vtQxL;�Q�v�����It�a���E;ڲ/\������0@�u�$x���J��Bk;G�3r}W��[��0ְe�R���Q��g�=�-+YO�³;Y�)�m�~��ǀ�F�R��0���3�V(�έ~�.O���l�(a�� �Q���>��a�����'æI�v����=���V�n�
��\�]%�ED]�����!��io:���^wlo�Q��|:&����c5;9�l�B�?��wj�0L]5��A�`	>�η���y�}�i�(��`gp�C�ѵ [!l�S�6���9{[�������^`�d���!�s�Mw�^�z$��4H�yA?>�dI"'H#z��a�?�[��������9P�U�͎�~{��`y�s���ᬀ���%�쟌aon��������ͦ�s�`�����f+Y�_��>�J&���B&��G�*!X���A|�$��ì��B�%�>?)�������`�:��!����bP�ĺ�ǃca>(ِ:� {�����,�Ԋ�ƻR^�����4a�jgۏ���$�]O�܏HІP�t�3[�x��F���u3���!@�''(��<���x�GA�VЌ�1���,������2�F1�B�Ab�t��������)�}��t�V�!
Q�W`�A҈�D����}ݛ��P���/���e�Bj�����~�C�2�A���x���I	^e"�Q��n 8�7Ǿ�ս�1�HiT�A�P�0�9ͅ������-4=��� ����!W�ʁ�6)#�d&��`~�(�uv >}ubs�����n�fw��*�a�fV��BP�E30_.��,�^+#E��9I�%�r5�)t������z�p���*}�z=>bN
���^��<���PG�dҡ�_�3P�xR&�_�F��\	���h#Q� ��F|�2v����-�4�O�xꁓ����]�]���B���.�!����Iu-I4��<��0o��j�o�-+��TG΀Q"9��8�����f��'����/�|WBw�m��c\�/�4�)o'�(�ӁsCH���"aH5W�Ъ�b.�)�d���ܔv�'%ŀ�|��v�'����	]<^���1
.Z����^0qe��m]��i[S+�Bj��z��B�~��Q�I��{|�T/C��&w���
��>2��s��yZ������V���A�l?s��PI��p*�X�o�
��o1}� ���!9��%��خ>�?�t��Ā#��alS��-S��Z��fN}�!��	�x�# i�����:=�F�!ߺ��:q\R��o�F���(�s �/�36�ٻ|��u��yb�˳�kii1M0�S�TBmzS�z���HW�]�#�2�`�&�:U����V0�c���	��_B�,��R�v{qהJ/����r��d�Jd�&4�vڱ�t�@��I;QE�s
p�8y@=Y/;����-Y�ΦvM6u:�ߞ�7��ץa��^�ץ����g�J��׺M2�K5:�#���DjM�x!KDBa���aw�?&�pm�FW	8p�,�|�K���1�q�c���� RA �c��Hf�z�EFx�cL;�'/�Jfh�aC:��?�	�s^�ʓ�Nuh6i��䗔�*3d
���f�L��;F�*���ZKU~؄X��+A�9kv��?�ܯ�/��Vn�2͚���s�})R.��{3/�]5<�R�&���(�84�4�[*s�D'��1�.s�`�#��@������Ȋ�Jm��C��1��  B�꬚Ϧ#Db~c��6���x�x��n	J^�H�{ܴu��&B)����#6F�c�1���̙d�W��i�Ք!7<�� �]^��qF�2�Y�6�by�P>�4j%b��"��
:w�++�+	@i�G�� ��Wi�̦_�c����N,�����,��T3]��A譊!�\1I܀vDM���D���mq�r���r��\
����;A��x�?z�?ٚQ#�3����7����;�3[
uK"c��2 OH#��ˑa�UhY^
�3D�� |�����i�=8k��~�=�`Ǥ
59&�ݺ܎�����<�J{�T�HlƧ���v,+_%�P�0؀c���~�A�p1��t�֠>�h�����Ch��F�[W�<�D&PePٸ�b1�%�ކ�X�E�
%45� �·�U��� ��� Ֆ�K���p��X4�cR�h�_�*��i��Nz��X���}h$CB�9�l��K!@h�eIk#��I<ޖ�)�0	�{&�s�G��B(�sE.�򅤼���%�jMM$�f9���\���݀!25�cY�վw�Ï��%+��fGa4�9����95{{e�w[]�?e*��)s�/AU�������R�WY%�9�be�a��~�Ȭ[��^_�<��h+0=*�TcCy�����?d\�--�0�սw��L�f}?�����4�y��myb��sS�`�݅7���5��<�dᶪ���rv�[�T�S�5��^k�W��>8�gb�8(AARM��+�w��A��P3e+�"�H�o@u��B�]Y"6�a#*��=�[캆����7���a�f��wS8p_Z�bTg��wԛUBF���� ��� v�J�ӣ�l0�QAr|۴<yڂ��|k�g��@�Tdy������C]�=Ӝ�>���;p�={���-�BGS��SUSn�v�ҷS��o�?R���G+�ga�"w�g0��h��B���j|�y9M`'ʤ���\~����g������5~xE��m�Q';	�Ř��w�	ܶ��G1d�ŉ��w@[�l@	�}��nౖ����
�|� �����&�c82=�'/�<���z	���j�h�u#"��t9��SD���Iꍤ��Jv�WW���{�Aӵ��,&��J��%��r.lRo��<����j�4�2J]��pή�A�+�	C��x��WQW�)���1g���XopE�/��ym�Q�l��R�]�b��:������*/�_	�K	�MR�}�8����'خ�6�k!{��/(��M�^镥-yhq|P�Lǉ���Ɋt}�Xq=���N�tT9�Nud�u�03\`~!sW��ހn�~$�,�z���%{�v�4ʅh�b;�Z�U���s�+��;-Oa�̐6�A>��v��?���rY<5��Oƿh��o���Z׉a`w+���/+D�����o����)%Bq
�pP���������25��4$�z8�����q}C��!�E����vYm	#[�����-QN�0��s���������P�t����
�f���ml"���L��D��HG(��Na�/���Tæx��G��!;Xph�/������w6#�Y�L(�P���aw'��'�	�qvui,�%f�A�}E��)�i�\�ܯm��q`�#�|nX���d {�5b�ՐBO�y��8�9O�y5*����p�8ld�n��-x��NU��I�?�2�EEs߯)
�7���NE�/��<����մ�t���3����p:@�+K�G��zE��z�1s4Z�!�D�@�߾�-m4�>U�	X������m%4�=�:s�Vi���"�Ǹ=��N&c���ic_�و,��nc���yk�;�U8F�z}��]|v��
���~���%������:�@���M���:Br�w�~+���޵=q��=;�s�&�y�[f:���gM�Z�2�ILYX��_����d��
�ә��rӤ�߶x 0HFMP\�1���Ъ4w�A�t�xTr�*�x����*��N
�F��X���m�s�#���K���饊��>UO-!k}ÿ��x��c���$폦v2'"I{���0b������[��Ԯ�g�G ��*��ۊ�܎���Q�ӯG�%ڛ��̝��V�s)�X�v4�e�O�,W�g$2K�+�r�&�.��0��_�lCR��3�)!B�x���fS�������W���䨫h�Z�l@τ7�3��l�<�@��'�A��q0&t�X�I!����SO,1%v�s�
-H�TS��R�!I�V���H���r��rv�!�-��t���b�zY���t	��c��y�8�RV8U��3��9��i �GE����r+�A�b��s����"��W ��7D�&��n����~��<��¡a�Ϧq�)�ӵ����K(��dPa����}�蛅��|��e����u
F�n�[�*��Pp�@IG�H=��<��W>���M�;i-Viz���L��5B߬:;�}�x�IV'P@c��~	%����"Y�Pb ���q��?R�U=��L���*�u�*dl����*���W^:8W^��.����o��}��Bef0ə���`(�&Y?%��R&�Źv��2�a��!N�E��\f�/��e�o�]��RE�m� N���0L5\�,h���!�]QA$XO��P��=C�n ��.uu�^!�:jRS�>@3�q:��	�Ԕ�v[�6Y�����B��D��,E(�=�e��׷�vi���	�aL�t��pn���Z/>�ȯ��he��ޖ����b'�"�
������Q��;AZ.�7�Q��mR�)�j��X�'4[�i�ٽ�@�ԌA��N)�������Y��R� (%�g�G�]�5V�g���LU��Y����豫S6�w>��៶�U�^C�z|�z��$o����Dl��7����.������9�*3�<�d��p��6ٗ`��A�'�u�+���� �ʩ�$�3�l(sc+�W�®g��֬y6(}���r��$A>����H@�q6z|!��h$Q�.t�ƊԔ���o�Z��+� ;��Ārؤ�{}[ �+g{a9�����`������'+Ou�r0g� �]+�I6���3(j�[�����󲑀�F>^�`����q�y��'�J�[�*����	�Xh�џ�M:᥷Ig�"I�龢�
T;�&����˩m?QHĬ��k�m[���!��M�D�i�h	�B�B��2�+����JƊ�_c��;�g���\Я^*�l|���B�H��!�9�Eo+���-3a�	qv+��X����Rq$�4��bS�v�AtU�߬H��Tĩ`z�l0��p{?gyz�S/�6��h0(�R�w�@��k-��RgK� �S��>���
nT��z���&�ٰ�Pɋ�~g�L��N�Wj#�N�H�e��n�������^�5�Y3_�+M;��}ʅ7^��k�}m����Cb0	%&��M��&�Ng��#l-1��
�����F���w���h�ė�+/�c�`QGe_��J;[�M���T%V�ߩh3;e��{�M`��ȋ<]�էKFJ�&�g�:I��j�AhEg����Ԙ�Oﴻ��=�C�*�!��&�x���{�5b&?�΁uG;��Syl��vQ[���vڙ�cl�N>��	����l�����5WWTV��\�[w�]Yw�6Bp� ��>м��md%i!��=��2�P����M�OVh�;���8�NGAļSG�T𓵤-7��9*��� <�M�2{��+��OH�].�*��%VZ^�wK���ȣ�����̽N"����$��֗�7�ť�8uD�1�8��eM[��JQװJ�5a<`!��&2��{#���v%��ǿ:���C.���q7i�+^8�4�
�D�$?il`s^�߇E-�qDc���^����q�K\�����N���������cu��(z~P�]�1JP8����W+D��k��c�e���4��� ȣS�
�nl=�;:��9�8��� �������V�Ry��XH.����gJ l�̲]֕΍e�`�C�/U_X6���i"�:�2�#�l )(�s��
�M*��B�<ߐ>3��t649u�E�}��V���f�e���QX&�]?����}N	G�z��ܺ��_�L{x ��7XoIT���TN'�2U�_톍sA�y�6/�5T(�
c�ݪb���Έ: �ӈ�,����e@[c�����5
�s��Z��Ƃ&�|3`��]��PT���u1����YA��?��-h�>�2&NI�)Lx��*�#�e���C�5
���*L��\V���ƍ���wC`�d�Os(����K6q�dĨ&N��2�%z�MO�Z��Ұ���Lި�Y5Ⱦw��kfh���%�x��XD�^|�"����
���MV�H�H�F\|����B��i��i\��7^o>���$e!I����&(��<K���p׎��%Yo�'<�A]֠��ba��=j�zL��R��[���.^؝�]����4V��ђ���Z���{�7��z�ʿ}_ۈ��*w�C0�;I+l���5/!�.�e08�.�]������L� ,yfi\�Q��a�f�lt�R$�AT�dd�����F�)���g�[b��8���VJD�T�K��) .�D��%U�DE�lE\������
T��d�:U��K�~ݸI(a���eJ٤�����!�@�WU9H������ߍ��ClN%Lt/�[�U�ᬋ ��Lc�+L��<z��D�5�!ydNq��j���t�m`�;Xfc�FY��b؊����(zl'�~���!��޺�C�:z�gT���$)�����^�	��T:��-�#��;�+ L�o��b��W"��]��i]eNG�e���
���X�S^y�|�O��3|���!���(��X4N��8��ǥ�ʽ�`��˟��S����U��y5p�-��0I��p���I���Q�q�" @�R������lF�%�ya�IX"�	��;��@�hY_�����;�!uAѪ0e]��n��eL�G���"�R�15f�Łv��<L�^������j�*˳p��z�G|{�G6C�nB�	��qM�D����>;�瞸+�V�<������piɳ��أ���M��PH�}Q@L����FH1	6x����f�R��W���E>)
eO���	��n�6oq���!�f�g��[��5��1��Dێw�"ƌʧ��m�ҿ��A��e� p[�g��
�ۄ�w��儯�٦|�x��k��cĖ۔������lg�n�U�s_ְ���f	D�e.%�o�i��%��|Bc6�*��[!��Q��,��
vZ��z^ڀW�-5�@���I�kO�� wͣ�<蹋�Z��"�ė>�A^����#IP��<��Z�yst ��.��+�F72\jO ����� 0Ӈ3�L� ss�P�c��o�%N�����0����	|�t��**�ŋ�˷:��i�04�-�`GN�� �c��I6��F�Ān��;�Ȍ��i�T򉟜�V�v��y��8��Mf�����vT�SK���"��ߍ��
;���xN�x��;��{������y&.G�͎t�R�lX��Z�(s<���*��qD6������?BYc�[b4�ʔ'���/�4�_��M̴d�Gt!��]B:�M�*���E��C�@��f2�6;̼0�aA��_+���r�ЦN�(6�bǧ'�����Ki���!��"�Ty6c^�f�ͷ*?L�x��΢w$npJ����Z*K��Σ��wml%��=+�"��ÇsBs���s��gir�+�i]%ca㟵Pݣ<��Z��TZ���j���Z�~/���Us6�UU<��8�ιh[�������~�<���v�8�k��$�����߫&�\ۃ-����T�S4�+v٧���#``��}\������~ ��
���4б�DNnTj���=:Fd�G��{h�w"��UL�ct��8�������C@&2��p&�<�-c&�휓��fO�]��\���&țde�C���<jΈ���,��ۨeN��Hj��������s����{wG���=���9O�&z���	c��t�H0��b�J|ϑ���������Ց��z�{�-~ ���2���h�K�Z*Q��ܿ�d�Dl;7��d��(A�)�?��7��5C}�aa�����:> �����|��O�jMI���o�B��k�\䙎kɿ՝n��Gq��݀���U
yC�\j6���(o�ꛜ�B�T�s��-���M��)xg�O����'�E�Qݰ�T��p�Y/��V:D:3���VP���=����Q[_9v�S���kٕv�n�r��X�we�V�S]�m��Vr�{G�`�S�j�yeO{0��{����#�r`�^�3f�)�W������/o�Չ�
���ۇN|��!eh0�y�6	��W�d�7���H��i	�;�0��s�ԛ�5�{��g's󦦰��3����SR�F��r�9>��bq�G}�t_�Z���V=+!+��� ����ㇷ��~����/\b�1pxቖ�*V�I���bf�|F�Ŵ!4.��}L4֎�䑴����|$����E����h8+4��0�̐ü*	�=XI1�7,.�*T |�х"^֪j�c�'�s �'����䆑.�
_9�z^�~֢v���1bk!�2$���6X�S;��;Wa<A�FG�#�l��9�q��}8��lDt!��PВ�vW�e��znW {C?4բ��k�z	偃/W2��7��jW\��+ �����p;�/����:/6�V���/oИ�.�����H��@��h��]?{:/�H�8���
����R�a|V��T� P���Ѩ���2�ڵɰ#���f?_���v|CH�_��dm$��L�kNK��� �7�s�U��=9��c�6����Ov�1L�f�v�?��b�`��βHp��"�Uڷ .h�s��z��&����8���zΪb4F�3���~�
���R �9&�L;k cH.�]k��FOQ��c�mS�B�����Mi�B C��e��R/��5�O�R77�Qu*�l+��(�����nd[�&�㇥&��H���+�����?8E@��]����R+��W�p�?�,������R��Hf��W��[�_A�<3��C�C�{t��A���
�;a�H�{1��j����Y�ν�ָ��z��,����7Av�0�
?��A�� �W���p ��f�Z9G+�\we{��kv�3�w�����;S8�R��,y��8O�_a�2j_')*�y�"pH{��]��q/��/v��=b/xw|��Xޏwj:i�պ��*�����_F:O���_6=��{DtT��xEl��"�q�9*��?u��4������ dx� �{�݅�l�R�#���N�B�ԑ@N��4�l��#W���I����0Ga?,#a��OS�N���
�K���޸��T#.8���#�Q_�H=�X�)<@�~�L'�x�͹R.�q�<�3ۖͰx!
Q����iD٢Y̨u*������9̞&��>&P!������J���Ã�1�
2�z_�|���P��������b�,�C4�Sը�e�o����p����|d������/��,�_���� h��dM��H��� ~�]SC���E)��M�Kmm���l�m�-�#�������12d4;�D{���	���u	;�{w�~�b]=��׿:�a��Cnj'\���ʤ���p���'�����X)z���ſ�ލ�
ہ{�X	9簄:U��'H�D�n��Y���8Ͱ2�M{��۪R7�B䖋�f�eDj3��l��&^�#hzʝ�2JvE�����v�o�����You�wt�2ӿ@�hi��	�J�;_�,�68���&�l���}:#�N�H�����^�v�U]5��UȤ	����(�.Y��0N�x�I��%�� �zU��*�vm3��
V�4��y��y?Քϕ͒Ţp�*eIC�~I�0�«(�'ӽ��OL� ����m<Y` �^Zm9�#��i�����c`����s�h�Rc'4@5ԧ}�p�*c�U��u��e������JO�֖���ewV,ԗ�ާyU����"����� |d�����q"���4򍑝�>(!`@�n�d��3�T畑ږ�:�F�����'�2���;������43Xx_[�^t/���>�4�17�ZPnj�q��u��p��,���U�7w��աӞ���'X��w���������y����<������Q 	�PEyytʣ���܆/=[_Љ0����N���I1ySˮ��(C�լ�y=����A�%�EʖV�%*�� x��M7��P/1��?��Ł��/�|S����8�ư\=�'�d��Us�h��ga�����+"��L	:���e�|KI�ݶ�]���o�d5�҈ٶ���s����	�>���9=1E����}�����vK74_?�1ob�L\�(ө���ׅ�0V���ŤdT8�ch�T���XpQx���sA�D�8)
C#U�!����29���5��U���6��}�!Q�4~�� �Q&�r؋�D�QD���^I<�_��nG̓+}�P\,ec�m�9�G��)>�/
���W�L�o����f��j�4��zԳʇW�v0p�R�{'�٫�"�@�l��V�2ԋG���ms�u,zPE�X9�B[/3�`���<W���,���^',��-R�2�>4�C���#�h]��U���P�����h����%S����]O��$�#�#y�;�!8�Q>f�\a5�97��Z�1��/�ج��0%����$o.�����j�aJ�
��$�.T;#/�oF�����;E�h{�6"�����צ��3�ˁ7Pվѕ�����_��$Y#��*��aD
�#�=�WR�xÊ��+�H��p8�B�v�3�	M��q��̵G��v�&j�D~���ٯ~|��x.;�Ю��aWd�zM���.�\i�-��:}]��Cn��������`������R����~fߞ\/j�KXˠ]l�^��M|��|�5iF�I~���K�mL�+-Ç���Ϧd�K��q�� 3�x��ɩ����C�.~(p�Eռ &�>�O���G8�~�`��TKn����9���h<}�u��
�5��_�H��+\8�O��f���������8�S�d�l��5��j;\DYgĂ��[�9�f�B�2 ,��̳X��өb�L��f/�O�U��ޚ��(�}E"	8׸*#�T+�����2����Czȁ��r���2^Z˼7坊��|m,C����B��!9a�r?ձ1`E����E��E��/�W���h�ۦW���%"0oU����/bKY5x0��D1�hr��֯��:2�����:�w���MB�W��3�6Q���+��he���ir1[)�!��$7��
�]P3�2�:D�������7���1v�hd[�xs�K|�S�b/�6D���&X�̑V�k��ċ�Ȁ���*'g��<
G``�Ζ^�@�h�*˩�mg����C�KR*C2VC���R�%	�<��2�:Y�-�����:��HR��54���H��?��=|�)άO�vS]�!#�ͦ��*I���7?44�aێ0�Fƌ�	����h,\*=�j��9���wL�#�!��ڥ%��;( Oߡ-��j|���n {MO�'��f�%�o��1�V�@p����+z������LF���I��`v2��·�X?��:�\�>�-� A����;�[�PgHYQ>1�5��o$�0Z*9JG�?��}�W��@:��)O~w��SĄ�1T^O��y�e��dg�@�nc�uDE(vZp��pG��"�l$z/:�"�~b�o"�'=���.Զ�������C��6k6t���Y��oo�˫��c�;��ZK�����D�9�5����Ͻ|Ŵf��Y�}<�>���a6��90)
2�ߘ��U����H�+��&��)�����^�ė�N1�L�y� jP��Lc�~jX�#�*���<��2�9�K#G�Q�Z���&^X�RE_q������W$�3%�sk��G�ԲӖ��s�]'ty��w�21�~�
��}���B͎����0I"���'�TU�W��ݩt,�8���BNc���;�ҥMug�C�[J��W���X j��#i�z�J�Ϻޞ����Tݛx��\�iP�ޯ�̵uA���mU�x�y�}�`4
9��Yդ���P\ܽ�WxX����ϼ#���E��E�q	y���7�^�d��;�m��!΀	5��4��H�� :�Xg�7x�m�ų�/n��#�|))�S�:��|�b�N�gX�t�&+/����˿r��`�I�`L:�m��� �r��Lm,"a�F}6�O�{A�
L>J=(t��V�+����N��-|&%���w�>�h`���J���maf���H��R�j(R�q��K��!��՗�u"���ɞ��@�2s%�J���dD�lRW�Û�W���F��{�M�0���ܷOQ#�x�F\�{T�G��$�5ӕ �y�h-c� �^�D��𳪩�e��(�b�gO�_&����6��ph��?C����(��ܻs/��,m$��O{��t�D�tX��/~��f�5;��M�t;�c��@;(VT�"a��@�w0[\N���:&���j�72��E����Y�4��s����8͸�(�1%6�&�f��Һ<��F���a3�Jh�㵛#�)���o;n�p��}�8�'ȱ�_s�D�')��
�rG�Q�?����oU�������x�'`�\ ��ֺ�m�|GP��唠�ަ��*�4�9ּ	��W�L|}��%��w���usz\"-,��%#��@��A���N�ƓL�	�4n=�ĕy�ü
Z#���=3x��2ԁO�T��q0��/{��.�� b
��G�ïY�ґ���&UM} '3�|[����oZ�@��.������ʹ��� 'iNt�P�Y�-�F����h��R���c�1*�`�,Z�e�݌v�d���PͶ��ۣI��%kZ!/q�}~�#�-�@T3�8�pĔ��EB'm�
����e�9��Ē�y�#�1>F�`��mv�=#&�n0Y�y���R�>m��j���ą�kƵ-�������/�o�ЬY5�.ճ�؀OSHS����BK6����O��Ok:� �D��+�g6wx�O�t�">��U)>/����v� �ӕ'�
F��"��7��_-��A��B�So�T���bSQ����'�x��9=m����D�"�iNS��N
ɐˤ��p�ޗ�?g;�Aq��u���r����Q������9����~'fY�a����2��yX��W�2�۽)�Ǎfig;<s��[W�����m��`˂��ӤA���|v�� �6�ܦ��ʹ#}�ݝb1��Q�����z�q������طGJ���c�g�!�H���ও�86�^�]}dF<\�3�9)���O�
�Bӯ�bU��-s�n���_����H˻��4��L�+�}�jS"��x%�� <��bB���T�?�(�u�#n��C���鶲~�!�&P��j�s�����&1#a�����j6���\�	�8hC���������_ý/��K=N��7oy�ۈo��e��'
�X�Ʌ��o��3ɃBe�;^�������Q��<A��C]Qq�3������l	�6���%S�y��wk�+a\	�V�p�*��.�0�crq@g������=��A����,F'�fp5����O��0��-H@�3�a���G�W�J��8�Rb����_ )���H�C��gFbxܱ���%V�˵����v�F�r�Q:��u�����tz-zVJÿ]~��x2繍�QoS���U> �ȅ��]ᘋ#3���2�J�q�/�e��8�_���Z6���aR�y�kH0r��2���@�r�xr�ԋ�eP���~'6m�gZ	alcYIu�ls�!
w�c���Ǉ�;r\���%N�:sr�+�x�@Mt�e�8�2eq��\P�D4M&sMl&��|qQ�%؏T����`��§�N�}��p;V���8�2���,�(f'@X��7.�~���3����Xc���"rD2j�[��[\倠 4(�i�D�K4�� �k}�+V�{������O������tM��}���������PLE�Å*c�ۧb͋y����ٱ�����Q,ڰ%���C��hη��<�rS��,�x[V_W��9�!0��uv�]�_viv�mC�\���ޜ��s�ϪW�-.�Aq`��xO�6�D"d�i<-}W����P��y/��&���,Y������b?�U��<�M��Hq��9�?�U������$�z�U����d�(u�H�@{Sop?E�A�����_6z�t� ;tXs.l�v�+սk�jѣ��j1gk�CWC��B���fR��$���b!�QR��/�k&sK;�`�4�!*u���Ʒ�}�?c�1s�E�(0�xM4�*;?9�cNw�Mf畀��|*�����;[�RЖt�׏]�tN?�ch5�W����v�V����Dg����W}���kW�YO�?��g����	�N�ؚ�!����+��Yv=�ws�Į1/�u��y��յL�D�h�=�9j�Ѩß���t��l���8����~Ed���������:�!z'��}�o2��;� �e����=�'�{&Z���=�(����ʻ~������A���y$�j@��'��,:qf�h��#�);MV)^x��/�$��*����a�9��g�
�zH���K;�D�:�[4�:�&z�lq��TX�A�`��X�%�8a�5z�Mw����GqE{F�2�G>�����n}�t�1y/t^�v�5l�ƟASa��M`�
ɞ9e`�j�!EI�n���懁o�*2"W�i��=4�uj��T�����x��/�4?<w6b�\��p\ø�("��rp�vk��)"�F��{ �y���¨���{vi"L`�V5���M�V##�B� ���&
&QdN���%�@)ˁ��Q \t&I^�y�/R�[z���y�@�R$�v�E��<ԅkN;���l��'
WK�Â�2n���	H(V>� N��p���=p���k�h��z�)�`�$��	J~|H�QS�� ���G������\#}&�[��\�- �:ۺb��<�3����g�L|ņ��G9H��uNMۃ�`��ץ�
�St�\1��`��ml|������*$�4VX�'-ws�f�~Sx�tZ ���*'�X� ������nR�a���F�-��]c7mi�?��l��׃�}�7%�.S[���HG��7j�fa����^CT`�$ǉ�6]C���,X3���g�A5:�E�\b�����]7����Mш{�Db���˾8��e��-���O<��%��q��G�w&v�Y��|�ݪ���x,�'{��*`N�"�8������.q"*��BM&��`)� . ��|H�=H�lc\}9�$J������m�2D.�W�5�juN�o��o)'��p�@���a
3է�7&�f9!�_�Ҷ�s�?���]�o�{@�}�r��<()ko:�bx}�gՍ�,��(�z[Ao��z=k���kc�Z�;�h#u�E)��`bu8�y�XY[�7��8-a@��V��g�Zu;"����mJ�h����}���|�?L��n���</p+��<?�P�eކ����Ώշ�WR��u���6�d� E� �*���\::jP��⠅d3w�嘉��&i�ׄe�
U_�p��Ԧt���(Fd\��֨Y�& �yզn�U�eS_�~Z.���f��UGc�>�/�����#��C�JFʺŤ�<R��E�-�2(����r�P{�y������v�W9$'}n�C���"�_�@R#/���r�W�;<3�QS���� 8��q���Ȳ���(M�Hpo�z![��'uo���?!qT\��UYU��f������7��.?[
�&0H�#6#R0�W��>y�FN�	�Rp�'��x.��������� �T�E��� n�Y�$�HX�M~S+��#i�+�)�̼�����]��27���D5�ԩ<{O adl��F�ݡ)3���^����D��׸M{!Q���!��/��g(�g��G���>eY��N������~Y�.`�W֬Ze�bI�&c9|�ܑY�~}��>j�sX*��~f���'��(P�ۅ�b@�?���M<=�`�>�M��_
�rS�t!�����=��7=���}�0�$%��r��~G�e���|m�9\r*�ǈ�� ޔU�ͪ)�q8�Zؖ-���~:��Y#t��a���:�ۊ<,nVE5a-W����E���1Q����v�G��jEs��H�r�p�*g��P��vc}!;B�|>WU����HW�1"P�\jD�>��h�þ,UL�*��g�+�����WZ���{�NV����M�%��~�2o���Q�4�oM�c%K����gF��Ϗ�_fU���ju�|��|�Q�l�%g��� ���Bf�8������'���
�&uձ�
�q�-<+H}p}������1�j�L1�˵��ʢ�	`�^�?��3dMa���i�q�@���Ʉj�9�*���D�D���潻��X�PsJ�dS}t�Lv/�bnm�_X�}�q&�B�Y�q��s�rvԬH�"�λK�?�-�fL�%�u+���j*�^���fV�I�2B3�w�CL^����E�_;�Z[��%-t�����Ц��*s�'l4��=�F�i���/�A�5������)���m�(㏷�dfDې�Tn�y��Tff�N2�K�i��$�_rE��������ˡRf�c\[�t����?�p��'��y䮍��u��;*K�"|�{7�j����w�m֋F=�k2�9i�y��AJ�;�? �� rz��G�]�TY6���n{=�a��\�3Sm�"Ak���uV�)P�(�����E]�������!�J5w��J�BPNi(qi�D,"��!��u���a�z���d8�Nek��
��O�5��OLN����)Tç�R>��R�77_ ��=�����y��s�V�M�}�ERB'�+h�?��iq	�y�@�j���ʚ���2�
�o;�;5�(ּٗ������jzC'��]"�I�%_	��M��Ae�\�����/Q�� �f��ä,�װ���EU��-Mn��l4�*�6©�7@�e�t�ƌM��T�NN^�{��`g�!�p(��z�/�{=`V�h����t�
��Z��eF�[C�z�_��]M�K*D��V�la4��<A��͈㘁�u��&-�*���Ss������]�r`�D���̗������5Ԓ�}&���= 1����oe�@5�ۘ�իu��k�S��XR1(�p0�^�1�}Q�W��5��p���k篋�TLL��������G	�lf��;VZ)��
���Ӣ��������Ԇ�A��(2��<���������7��1���1�������la@C-
��!Dٷ|��IM�Zut�a�{)DkU�u���Z�jM�����m��A���o��54^w�?(j�m�?�����ڣnEY����hfq2���Oa��#��7�)�4��I���T����_�Zj �E���*1��l��V�gt��]�y+h�TJl�����ÞP	���h��Λ#;{�Ԯt@�/���,z�wݹ ��C��]�^�g�/sD^V9��w�=��	q�Ji��	w��An����򱡀͘qT?�Ja_ u����df�J�l��v�7�F����,HzD�~-�;���u�F�G��<�붊��gR�3�AҐ�} ˑI���k6��*���BL2z �I��@��s:v��?�B4u��9��s඼@�c�rPռ�+%V�Ɂ�<h�C�s�oUqr���c3���	��+=��J*ꈉ�T0e
3C#u�h`�,�AV�qCp�/e©���~�n˜�Цs�X�26�3Q�:�����s9�1�A(�)�Qk�an����h0�u֖�8��qc����M7qC���2�'����;o;�c�}-����D���Jlq\�\�_��'��v�}CrG����w)V�[�j��C�/|�h�5���?��
����Rv��Q��)�������=)�E��{<z�^́= 0��.�n��WTQ7�	N�[ Hb!�F!Q�h� ���F8Ց�s@��M���$"��-5�-�c�(q�����(�5�o��R �W�Ԫ�����v�=G]V�""Vmö3bSxp��4Fz$��U�c�3�W�{Ϛ��x�;8h��5�Zod?���ԫ>�g�6\R;�'�����X�<\:�B#�'�ݐpG��h�!����5����%����85�Uh2#����~���am>�"</w�X3*�6|���M�%%�;��2>���e���o�[���$.ݗ�ˠ���L7Ü#�5<W��'
� 
��&��=���E������4�7@p㇔I�����c��Ra ��"�����/��I�gȤ<d�YXD�b������Ë4 l�\-O���������R,��s�3xt0��e�Co���J[���Y�jF�R|5���zX�+ª��*���!s.e콑���a�nd꿝uvĞ�j9�A�����v��^�/]�|s/mf-�-x+�]P4���<���gF=��Ji[��y��O%RW��O#k�8l�9*�?��w�31	��{��^[�7Pdr�D���b�������_&�����)N�^'v�Z|jx�ű@��o�y�%�u�t�M�|�8¼$ry�3��'ʪv�v��2'��'�B�I�sm��� �zBt}ƷU'���/�Q/r�����j��� ���[b�������@_hA"�}��f�*�7^���_&�8����Ҿ��@]�צ��FL]�b�� Ec��&�C����orN�rJ
�ڱ�(�|�pT���$٧�3��v~�NV���?�j�DAɌ�q'&7LY�U^�����vx�=���μiԝ�/�X��FVH��*v(
4�57W/6�Q���U8��V&�vJ:����	�5�Ӱ	|A�5���Z�����,�G(dc�7�=<�~>�M|���G��`l�<��(��(=0h�8�X�,�,y`9���̽�?�U����A��ڼ�r~(X�I�Z�$��`�?�e&��&:[݀�^��}
,�-(������Va6w��2��W�p�A�7.���{J�ʕ\uã����&�����ٝ.-?�oP���E�5���yekO?/�Y�+p0َ���,0�wLrF`Y��(��1��9�~Vۙ�+Td���K��)Q)Y~�ه+"s����.K��^�����t����d<W5�n��M�e���j� �u�
J�w��g'��}�3����/F���@��1�#��ޜ�X�U�e	��$3*�6��m�x��7�?C��8�<�,�/'�����9��i>��d��F�f�\��
�pC���5�q����[W�/N2 f6��;�)Jq�1l0�
F���q��І\vO�����F\<]�k��v��ȷ�\:a1�3�ɡ��@.��?K���uWo������ii�<���v����`7��o�⳹}'�O$��D���� �>� �J���r�y\@a�­*�f��4�j���s�]
��u��=�����}I��T�dϟ}�QH�FW�3驈�k[�v5��T��^K�]`z���aQ�#�� ''8-ґ%cϝ����rr6�IȲ��3���|���[�r�OP}�y���h��5�̍�0���H�jJ�O�l�#�/��d�ۏ_ebS��nL�5 (>;�E��A���I�}��t����x�N��T� E�"��^'{%��q��O���K�wZ!m���,n`��@)~y�!�]�����/�b����Y͟��6ܥ4_{]u}ᩅt���0sʃt(�M+%���Jۂ3�N�S���T2j6�{Ej:z}�	��sOG}�Nps\�0�z��0Nyw�d$�,��ՆL�|fY���������bh��X�"9ΐ�V	̀���e��p�Kf�g|�Vj�0X-�r�}�KK��sh0�[���+�;/�RJ������,G#?��J�0�7q����spa��rW���Rsp�I�e��y��h{@ŷ�׊l���4X3��ETsL���bV��	�� v��m���*�%�v���q7�������y�j�H���|�>�����d���UȚ�5C�Ϩ]��N�QJj�~V��K��ܯ6�H-N���Ei��*���g����3���l3�c��T�F�t������@��f�)iV�y��t\
\v��&�q �K�����H&"o�3E���X��w�j�8K.o�ةH��&
"j5Z�!G���:�_V�c��Y�d�%�$�u���O�3">��c��}����Q0I?���X�4�n��ip������uN@��OY��g7\�^ǿͷ�u���n{gp����kʐ�T{�����Ø.;��/p^Ԭ�����k꣐��0�;���Y���L�4f��ɚ�x�Ɯ�"�٪��7px���ms�ܦ�d�s�	�׼`�zÏ�����FB4�!(��Ar��V jvR�<��N�V+1��.IT���ve�&�̶�n�4W��%v)��E<X�%�$��m���4~�����R�[��T�|K�A�mD'M�z�]��g��:�^%9��#��cd@dJ[[k��@kp?Λ���}ƪ��F5�*��N23�"=C�w�5}�R�!��kC�
��Lu���^Gl�M�X���=��y��n��H�~j���$X ���ܺjKN�BxS��7���쁚��lB���EU�3�c�h�J��=+��Ӵ��]W!Ҙh�H�O> +T,`n#� l`��K$ӗ�e�F��2���E��E��N/g���Q䨽 x����Snō�$ϮN���2��s1ݩР��e�̝ӂ�:-sg%iC���#�Pt�F?f�/w��z	vf�[�H�d2��7�u�F�k��p�"���:�Vd�ρ��x;�%���r�S�5�j�b�c��r:��o��@�SA��E��4���b/�C�RF������lf���uГEs������J���F��܉�eL��<Q��>U!4����)�)t~�E��`�P�]A�i�p��=_<��	 S
DHư��f������ ϜcxwM��$y�$���>~]{�?���4�R~ L"���0 �	��2([�+������4L�C��fݸ<�⼣x s�`a���w͔�n�xF��=��A����q����@p�9&I*�w�F&��@�ǹ�AV�r�׌DT�Xȃe��x��ގl����1o��[��l@;�Ho'�	�c���wvz�.���7E�ئ̫��)P�;��^P��2G7Q9��Ȗ�#>׸�;C�V�׃��[�Q�<ȠR�/]vH��)5()#�t/k��B����� 
ʪ����.��v�;u�o:��5X�t���	�FG�]�����ud1ֈ�"5���yV���d�����H2�$w9��;8�#�k��5vs&s���l�fAv�nu��Ú�x�=O�U2N:���̡c��#D�7��n��|�����ԳR�q���k��%G�:̞2��Ft*������yy����_xy��zL4A;{c=&��&�Ke
fH9낤 E8�j�-�/=�p�,����ţ-U��CFف���p�F �_���VB����K����M�����MJ��O�~��x^���0��8��fٹOj� �K�1�y��j�Q�.A.��Q�
��;��` M^�H�V�e��	��.��S�z��R%�讯�
��ַ�:�guki�j��bs��$)���L����ӫ~��-|[,��P�%��'���g)��Gu>V�"P��|�}���)؝m��|��<�J.�7�z��Fi8dO �=������W�F� ��01_�V��<�L���: �y�,%�[�I�a�{����޶ui�,>����l�p^
�4¤���O6�ʽc~lc�m��K&�,s�$�
\6��Zw�|��
Ê����١�҇��Y�B,R��	>a�s�a�$a4WK�c�qB:����n�g"�]�af��u�k�X�u[o� fp�I��G(b��/�I�����U�.�Xr��hH
H�`�nOq��8U���ú��o,[�fq�/�A��$�hں�?�	��c{[h�`�Ao�]�U�����.+]�52�NBD����ʰq�W]"�^�C����y��q�0b2�k�f+4乐�r��W�gڡJ�$q������@p�[J�Z�xW7e��A��1?R
��S����Q$Q��'7	4 �5)�Ǿp�"�i�Q��3I��Jp$���6J���	�͹�ֲ��!��Ɂ�U"�t���g�������iTۆN���z�T�r���ޙ��.Ḍ���G��.�-�����W�_@x�np�dGV��t�M�,�W�~����5�툫`��Iݶ��&�=�]ˍ�Vӽ�3پ]Pm��#��z�������op��˰�c�׷�j����W�q��ܙc}DA�a�Cƺ������x���OI�/qb�U�s!�e<.2lB.a h��*V�� N����K�k��Oʭ�͟y%_�����R9l�z�DV3��_�q+|�
�ȱ	�ؠ��@���v9��ed�U ;AL�O[e�4 �g�07�������w��2�(�ټ�]\�RX:]�'�Ռ�������O�t����PG!wH^��ւݍ�x�=��6pXw%P�!iĕN����}u���Y�蟷��"�aTبE�w��i�~���:Z���H	=��}�=M�+;�J%1M�]3<����皚Z��ч��I�$MHRh�b0]��ֺ<*�#�Z��sc�]Yvh�����6�ԍ�����9`2,���	�Fy�S�$1s�?����u�央�-O���_�}M��}��m�"��t6p*W�bI�7�#��r�
R�+���m���j:T��bd�ږ��� �.��{ ���=��n�Q1�<`��P�����Fn6�8�b�r��d�)*�/J�>Թ˴�=��|��3�ea�c�F�����H��^�����C��3-i��,#�Ep���HBgO\`���c���Wh�wn	n�r�D8���_�y����Π�G�,T��Q���y��~u��N�� 
&�����$׭>�$�O���㍼h�2��0O��f�LMw��R_�?Yw5?�0���i��W�v���":Wt�5�;y
0�a�ę���zvD��ZcX�".Y���2$����}I�;���6����㬆C�M����Ǎ�-A�X}�<�4M�u�h<U�S-O����3<�=W-��н鉽Qxl�>�J��r�M3��l�{ռ��
�G|.��>J������@v��c�r��A�'&�`��Z	������:ψ�����-�|��?~�׊�����}Q��	��zA�$���'�$^��V,/fT���њ3AG��z|d��v�k�'�U�G�M��Kr��4'�h>@NcD�f��W È�V N�)H��	�\"�&˻S��a����%�����4�����}c�i�#�Жr�#��W�V4ʧ�3���Z�h�{�QTWM�?��<���nM�_��^1�`ڭ��#>M��&�F$}�o~�r} �{u���&�6Ҡβ��_�R�h�0�l�N�d\9E��A2Ž�����+#5�i�����A^���7�05��E�Z�7	�N��py)9-X�"ʂU�U���A���&p�`�������S�`���������~H=�jҮ�,f�8(
��2E!��Tnv1�P���r�S�Ϙ)Znh9��O�G���w��T	����y���7�9\�oug�N71H��Otڄ�Pw@x��{a|Oj%h������;3w:�|�S���D�!���&�`>{��Lz ��g�r�X\��S[8^H���q/.=Rۏ��f�K�G7������g�Y�L
i)qo�6[��w�-Rm�+�)Sj������`�+��z0F^/^�K��S���]�S�>�F���� %����T<*�0a�$�4�2�f�H���h�C�*�b8��Ĩ0��v`��u�N�;��"�=����9��H���CѮK-�
ڱ�o�f	����Bp`P�,�n8���0����_�`Ş�3B�pۗ�nU�o�E|y��׽'iսRy��<[۠ɟ�oS6���p�>��!���se�8��7��,c�!�������̀����ο�e���@��(NL���nĒ��B��SwnE�r�b{� ���}��IB[�`�Tt�v���ra򋜱�Ol������܆�1����vG,(��m�|-��j�h�C�oU�&"w\:]�}��ٍ�Eam�	����m�����܄��K����W˻�Ǯh�E��g��JeŞ�C�M�����T�y�o��z�����1b ��$
� ���W���&�L�y\,djH���m��r�Ǡ{�����7��K[�	'X-�cJ%��;^d�j�f�@m�� -=Z��~����:}wwgX4����%��@�F>☷bF��s�Uis3���,�Uo]��ōR9#x���H�IN��Ǵg2I3c�r� �$)e�͡O]�@]�f�M$�_:6I�,���atR�Q�=���ۓ��cE?}�]h�1�F�� :�tl�O�?n|\��C�$���BpF��P�� P̻�^��p���=	�ꂪ�ޮ(�}��S~��Yx|��eQ�G�E��PA��
�!��p�m�Bj���"ؚU"�gT�^ʰ���� ���¦	��ʚ5�y�#c[�P��8<����:�1�P�O�;}�(1����t|�T�ג| MZ����&��i�l�h�o�s��Ovb�d���4�>�QDQ"$$��&�9mvF��ꘊ�mV�ͱt�c�(�ǽ��n��`tͪ�L�֍��;�=�Q�����miOlTM/ ? �ԉ۴�]�k�
�O�N���e[u��b�a/f�2���*��iK�I-�vYh3��F�X����{��m{fu+!_ ���&��me� ��dT{���FY;�dZS��3��nZ�Qȧc03@�z�C����7��&	��ܸؕ��FK�"]U�� s��q��^v��s@<�O���hS��N���e�ӗJ s��h�1֚�'�\����@�Ix�x"_����]��Js���2��Of3*@	�3Pv��V��11-���M�8���/�!JCs8@�#@��3��v:Q�ӈ��*O��=�݈T,/I�܇�N[�gw�EPx��%�Q#kKo��x����_NQ=�M0�@���x�Sn��܂f�!vT����&a:��>!Zd-T�͝es�E�&t��q�ؽ���c�B�M���W��.߄m-�f����5���������0��hp
j>�↶!n@n����`���@B]\�&h��O���<A��fI)I�:��-�S�2��vc�Kel�F
�_�����j����\�2�ܐ�����,�!2청J�~��P�m��[�2٨qH����od��4�5+�%��'N;"iP?V]���a���I���d��ယ�S��ΚB��	pH3��Y�����l��_���b�/J�p�t^/�����	������E��E�`"}V�)S�fê��2��LŸT���s����c"��wRBS����a�+���h����!�wk@���� �F%�l%���ڹy0�(ͧq"����#�m��h쇇�X:.�za=��З����$.[�0���=k�P`U���O($�[,�M�(#���ou�d&b���R�"�;��e[��szs��Pb���� rm�@��>.����?��Ċn>he2�ѩ�@�<���]��H��w�yH'����龈~P��/Na@Ԭ��-i�Q~��݉�6h�e-���l؈]��DX��`u���S(�WH��G��Y���L�����N�.��|���< ��f$5��s3����I�k�k��i{���@�G�RsAJ���&+��t�ߡX$�{9K�TPv��.'�}$gM��ћXb)��{6�����y���y+I4+O=�l�S��t�N��z��c���{*u�����d,�Potx��=�TЍ¬s�iKJ�0������(��7u؄�)H~;mV��N�u� �Z��N&�	�@KUE��}�L�ߪ+�O�k�a���[��A��:[I?A���pP��"���W�F��Xg݇4���-V3n�US.�6�愼�v�e �Y�]|��� ?�6/���4�(hS����Y])8���>�{��q܃�[���V`��7o/�S�n��+-(ʭ[�n5��n�W�"�wi�tri�d���@�V�����׬ �F>��'p���_�h-7�o��S����f��Ͽ�rZ=�Zt�	d��S-A�6^�ANO�j�����G�0ac�Pv�a��y�p-�c��_����%�r��oK���{%YԶ�޺C�C]i.+P���~�\����
@d;x��t*��/l�������I�
�Bآ8ש�K|N4�֙&�)	�dv�__� D�`(uW�$?ì5o�W��튉b;�%-�W4�<?u�)vy��2x�=:���m�'Y���j�u��S�R��h�����V�9�}CǸ���Î�_*#:�ng�yؙ�Yԓ�>s� )����c�e�?%<5�� �q���Nqd��$��d�$qQ�
>%��$L/l���^�KC��Ā�����xMA	�/�(/�QD�� [7[��`.r^Ұ��Tx)��Xx~අT�bI����;���WlVi�Vdm��"��8� ��,uE��=�}1
cknUX�<�O֫�������� &��t�x���0�eOھ1����a�C�����%���J�Y R]��0�����*��7�+^/ s�^�LO�7l	$W;����E�`�OяiJ�k(�-t�֍5�q�t��/�K2��*�%7�!�y�0�2����k��L����km�p�/�����!��{G �\Ý���ҔF�����	r�Y�mL�<,N�=)$�Ir�Ԋ71<%V�N��6<TzOM�5Som�b�a�@��HQ�+��-9�/��X���9}߫Rx��1��l`��ܸg2n?(�7�����i�����h-��n�t�Q��;	��ݥ��S�E��	�S7
�w���5���	n��I��A��_
�������P �Ѐ]��Bȑ���귎k����4��m�#;�=",��2��i$ժZ[�G�ȫ�)N(�6�B�H��G�WyV�� �+"�EB�S��m�DS������;d���u����lQ��S���;�sL��K�$�{�}�D��w��o~$�������LJ-^r�=T}p�����-t�"(5�#�%J��^s�}�F�'�`V��jȧ���[׶vWؗ���X��.\0:{�5�
�<Z�o���WC7�X~.��& �j.�#��M:aY�y�B"��^�ح6�5��Q��;e��6�"�py���ǯ
v��a7�]@�V�B���	 �?#�_!��~���%&
-1ᖼ�ɐ+ȢI��Y�Ǐ�d�;��^�!��S���,��n��z��[��o?E
Y����P��/���<�$`P*�㷶4�Ǥ�|Վrl�~��7��zx�U1Y�n:��&�<hdX�]��צ�r��h\�\�#<)x&�[�� ���	��RI�ڥ4"X����d�3'������+|������~br�!7(�`�|ixᶀ�3y�7m�Xr|R�^Y��3{�Up;F0�`�\�o�)){6�X��yT1��39J����Q���Z/�8�=��_&��~ܻ��z}O��T����m���d3YeХ��l�?Pn�fr�ݬD�E��3�%��=��6xcf��ۘή�;(3�&=��Mm�O���.��\.0NS��Vh1�{�_ޗ�|�w"o�<���7��~�xm=��,X�f+h��S%N�����χs�Շ���!2I˫��C!���^J+D�Dun��ǽ�DwR�jv�p4�
��}���5���KN\�)f!���E��������h.�t����Bn"�06���tjv� �\��_�:���ɼ�Mnc�/KKgb��\*�`����؛��\T��5��ݖ���`y�	@�a
��kV�9�������U�\1�$�s�M�G�6��y��6�J���W�Aۘ\(H��Q�k\Ź9��86]�\��I�N=**^�:s �F��Fn��&F����S��>���!��='m'�u�Hĵ󶝮u�A��H
�˛w\zv��:x)���'��Z�B.��	���p��j��x����vkD����/���&!��:��>���$'�v�{5{huA����Φ��E2a"�g4ݦ���Txy����?� ��l����_��2&W���
�����,���y�<B
:�qip�
3&	Z�0Af� N{|��ɼ]p�*	�жP/z�-�M8�l�A0���ς��'��-B1�Eem��{̃�#7���ߎ?#�ed�2ɧ���q��Y�U�`'H�n�2Gaj�2\6��!{�zw��^�,F9XZ��a]�2;Py��f;�������t��JѴ����em�/ts�κ��K���f5:Di�:��X2b���}@0S!�ZУr8�騤$�)�H4x�9)���'��J��Pc��2�{'��������E+�{��Bۦ+4�>����M��gt�-]<�?����پL| �-�0���:;�Ͱ��l����|n�l�f����1��⾄	�9�8��%o��ߠ��7����h6j����0`��==�X��)�4���,�����+�FṘ&���D;��I�8(7N��Z�j����<M���/ ���e)�4�l��ts��1F�G}}[�BQ�K�����4�j�X~|?B�6�|����� ��3��t������s����1�E�#�F��aۡ��/B:j�V��f�\�?�ȭ�a�%Qu�5}i��d!܍͝3:�!su�Y/�=�F~��j�Y׸P��Z�FQ�Z������'mT�8>6��n�,Hm���r^ް�����h~��'
D׊.�v��>�F���T������J���:�o��	��'�����/��o�*L������
	��&��1`H���<���k�d������{-g���j��m�*��%L@ƭ;��df���k5�I����X?�W��������Kͪ������������_�k��9h���Tl�jx4��r׭�����pط@v�-�����tn~���*D-���g^�D8 H9�4�g��r-��M���MS�p���%����t&�� 
(�F� ��{��_��Ҏ���ү]��Q˫5�\l��c�,&�Wl���z<�c�POC���F�策�A�b��H3᢫. ��{9���W!1w(Ǫ@Ç��Y��z�W�\�۞�쮎k�f�i 5�λ�XE��ŗ�}"7ݘ`ݭ��F��"��qG��;��{;��L�af�~"cs���I�s�p�ǉ�\;��2ڤ�����GF�aO�=��^��e�`�
�U�2�!��:m��R��Y�R�������< 仄hyW8<{����c��N��z����gI�<��@�]H�"�����<�:�k��*�lN��dR���q�9���q�_�����W�a�'pX^�����+0��F8jg���2�`�����OQ�I�ԉ���E��a�J��0&Di�V����p�F��t(�<N;�](S6��
/댼#�����s����/u_� ��A嵼���y�9��F���|Q��c�!_�-Y_�l߼�X�_�[nM5ͮ���,jq��+������S&!Q�Mh���ws��x]U�'k@�s��G	�"��zC�gU������� �704K4���&B����/�����8�t���;_�\���Q�TQ����ȮO&��h}�%�yj����}�Z�b��i���xnW�V�]��3(`�W���MF�(x�]�N-(|�Dܳ��ӓ��$п0o��aSC-�w�F���5��˫�O�Zv7g���n�j�yY�q	����Ԑ�/�A�gst����C1�V9��!y�5�t�~kv- 	�j�=��4��nGu�<98���YD�Rz�UsE��Z�K���bQ6gyF��0F'����>�S���9��?R��.��C�����j��v=�M��-\~9?Hnn<�LyJ_"r��ï��J���K��M��Qm���*qc���1e��|��ɺ���S�lg
���3y�cv��9����ժw^��k��4�k�0� y��+|�ĝL��oy��*H)RX�
���Q�O� Ԝ��L�c~��Ghk�K�x��a��#�I.�,�h��kR5v�>�_����������P%?�d�<�V�j����?��BR����Ҝ�2��*c	:�)㔚��f"-��H���W�|&���}��� �'�[�"��
��?S���[�e
o�>�Dew������iA�#�3k���_�^���eϢ?�aG )Mf����b����F��Kt�1����rC�=V�=�/�h;<g	�3I=����Q伤}�I��R���]�C�.F���������Ooh�M'���`"r��#���m�g@��Ah����0��͆�ӂ�F��yy���^sK1���~����%%�P�����N��\ٮ�X��\}��s> ��q��3�lkL>����d17d��ȕ$��ì���� !��w`��5��h�ϰ�5�DGpw��
�$�Y$A��H��(N��q. �������-��u�^��+�N����3x��sg]>��g��l�O�m	��CW0Xw���𜌜�%~i~��\�{1V#����5#>D�N�n�}vC9B� G%\�L!g�X6
�b'i�0����1D惓�J�M�[Op���V�����WɆc��T�<A2?R��[��V�'sZOb��mX������(��y,����l��Sҳ�Q�Qm��F'*�IۉԶLʋ~�����p�i�e�U��a�W��2D��ۘ%�O�9��|Z�j�(�H͂w#%��\���-/`W]*ͷ���b��h�,e�Z�%����l��	��8�������?�<-��o_y1 g�/�G�n�HU����	/��k9/���7���	λҎ�JS�Sa�d鱍T���m����b�a�_t��!g�[���L٠�đh!��=z����y>Z��=׋'��,�g<Y����)�9F���ԟG,��,��i!H���2iu�ֵG|�a #6����9a���2��s�+��J���P��/}l�a[G�T@��`��o�u��|5ZL����>�ȉ*q�hQn�L�Vg���7E�{�v"{�4 ����1��lC��e��C��!�	��o�ν�%���/�]���vw���)�ւ_�MB"����LJ�F��Xԏ�	��t��� �?'$_��v����M⁅��7��8ה��ͽ�D�_�$E�dF߹㜜c�T������C���58���P��Ĥ���)�D;�xS& ���e���H�v��
�,z�)��2cT�%�`)�XuAW_J�	S}Gޞ�/T����}�8�p��B5UA�����[�e6�U�uB��H�����*B��^N�g��{�;&�I����@f��Aq����j=-��H�
EY�Z�JF�NZmNO�
{���N��7��k}���ϓ�,�|�̄���4*�x�A܆] E�F�{�>�Z��ZZ�Q��|�ni%���"�V�>^r?����Т(���H�qS+Z���62�`�Q��Q�Y�d;X眻`%�eO�G�0�[ˋKKУ#U� �2�~H�U����oߥ�"%>�e�d�NopRjMu'Z��h���=Yd;xt��RI����O�s�Ϛ�G�W��n�t��O��!rڲ��딧Uڝ�p��ݢ��~Xq�ݘ�b��9����zҡgU�3�'k�0eF���!���QޕIiDsܛW���l�g;�Ս�Hr��:�zvL�0y1ʅ��ui�C����lmu�N��{`�wF�_I���a1��+@`��=x��fQ�eN&.鉿�[�5N�6� @��c��03�tfÿ��L�Gh�m8���{�H���v���iѻ��뚉�9���}��_�G�-��4�~j�q�� �I@����nz��U?�5�=��s���N��n}����b��~:�;��{������7�)��|y��ڴT �$6�5���O��6����3!>\�o̶i���.�[��J�܏���7���NѬ�,T,�kƕ1���<����t�]�J��tu�np%�Ě�\��4b̶?ͼ7=d���?���'������Z �[� (�L��KC�}�Wk����Q`u!��-��k�i�E�rd Қ�&a����1�.��
�sR|᪆��Vx2tJ����mp��ո���ʋ?�o=��<���g"vr�ȭ�1.Nϝq-�(����ʍ�e�g�G����|D�$R�&W�X���H����������8���$�.���:B
&��D<ZU�.af�[eG޾��hC������>��a��7�wU��;��/�~�ls`?i�Wh�[���L��Y��j���Ý#}U�b����pi�����°�BL�3S�e�35.�l��[F;7^о��h���)�� ��8˿����R[@�]�_�]�g�T猪6���� �1�6�)4�Y4㾍�R)���<p�Eb�j�ЃD�AJ��+�!��f�`�)Ʈ�V2�L�<�ǅ��ax1�k�$3�g�D��e��eh� �!�<LFR�8$�Hj����2����aI�-:ܻ�0��Yڲ>^�����H�.���O/�!���jpw�MV&�ᛊh��}P	/��9��!@\�\���B���J��ȧM�{�[�/Twn3v
=䪘m)Uo+�Ŏhւ[z�YR<�s�$ߋ}�A�? b�S(���QOe��aH��HPn�����JwI�a768tt�ؠ#c�/ӳ�'���z �(��= ��~H� ��D|�(W�\�\'<g�U#�8yR�4O�8�M�I�p=���0D��;(e�.�e��0��e �<Q����"[f9���Z����J2�����S��m ��"M�d4I��b����FlGM� C���-�]�a�Sy1���O���J��g�ա�3p�S�8-��p�oQr���_w�Y=��7��1��o�'�Eo�VE;ó�P!���X�d�NҖ`�R��2�P��v仿�U����mbH�Z�jޞNajKF�d(�Jm�C�[�z�#�5�g���
B@"�n~�c�)��$�1���3rNg��T}�l�A5ι��"�?#Q�Q+9��_nA6Cn̤*ofN��m�8�S��94�;�Kd�"אY˲a�5��f�q�n�� TE�c�d� s�Y2��Է�0�]���v[�	�b	�_��G��+L��0O�o~-T��{͹a���
��U'��64�È����{�l�ƹ��a��ߍ&ú|9US����b����'��~���\�<�V��qXM�`�k*2\����x��>�����]q��B|P<
/�53#�7��hsk�d���)�?��!�wr���}�:���G ���CȆ#���n�_ad�'�JS�*�U	}k^Bc
$��NfD��vXV�QR���\�?گ ��R�ޒ��N���Dz)�*EU�\QZ!�&Ѩ�!�s~t�����
����
��b(鉄���ȗ�����W﹁`�:�w�Rw��3��b/L`ғ��)Z�г$Ƚ��J�TG���Ӄ#g��>�И�c0�̭{b���_4!A�Ƅ�2Y �+���|GkU�OA�sO��Z�n�ﵱ^���̣9�����c��k�F���8?I&�$B�У�b�G�4����5�k%���r�K�@��'�Ġ�
��l�?���Ui���(렏l��uXR˱��mxB�BaouV�:���� aĔ�ew�oI$.�kj�}F����KI����&ܳ��Ӑ���Ѹ��9v/pB�Rp���z3�
~�� y�h��a%��GҮ
R����u��7�Yl���xI|�����f!~��A8�k�O��m	Q���G���З�~%��9�w��P�uR`���=�ut�W��0t���c��T�����@R���
{��9
:��g���/�\S��Ҹ�ri�.V���!�)�ѷT�J�G�jk? 2z����D���:��mrL`m��d����(�������c䏁�O�S�6�+��(����Z�Ђ�6�[���H��:��X�'����h��S�d��m�^�d_�'��/��[j���͕8�VZ��5����d&*�y��똳mf֒F,T��%��ˣ ���D�m5�d�9~�o���NtB|28�N���v�8�,`��r�^����7���,��R'�U�-�r�x�ْ��&Q^vm��p�J�a��&<1�:%B�@b1Γ%+u!�Dީ��mBY��d7�����%}��d����s� χ�.➑��%�gh�M��[
wX4�X�Z�M�V �*�6��"�t:�-a�`�����z*r�<u}��V"����n�٧�͐h0�s�W=tb��b����B^K��]H�
ҽ@_��O},�fSz|�9n�%?�[P�-��(�&'�e�hG3�&gX��&J� ��R�Ċ2���]4 >�!��6'�&�v�;�p�e��[��:U���1�F�sy���W|��@zU�3팖�2v�e0ނGW���"}K��.���wd�u��ʸ���wPXA�Й������9Y�.t=e8��P���N�6I.rp�4�Zt�ve�LO�rEh�G[KbZ1J)�����2�|����Xfl�I�[JO���$�N8I�^�����C�K0m�՝��/<� �M�,�d`Cc��p�(6_�4 ���\��? F�ӫ5�3���9X*��O�;�Y)�?�9Ʉ���ױ'���*S��v��̖���|�EFL}t���� ����%�����N�h�����.��<�Y��CN	?������N}���M����&��4�+L�}�a�bg��ᷩ�`@� Ѝ���@��	moA=���/#�gW�^�6������!�§iNs�&z���4�`oq}�l`��&>��;���A�8+'�:A�;�	q�:��Z�
�+��?}��Ӽ�\`~���)�H��b*ԗ$¡sY�*����X�\-����V�׳d�۝������q9�w��b���~'���(�T?zG�\u��/�I�����{a�J��� �	3��mʱ�\�5 ��j�~{���	�w$��m)�V�v�8Q"8�ĊRP{A�[~x.O�˦�JL	�pAI��K�������)L�E�f5�� �]�=����װ�?�C�OBLd+�y&D�1Bz�mS�2^�J�m����9��x���{6�z&_*�W�D�|�i3{G��g�{��RŏX�|��@E�V����;L
��X�ͺV��u�5�����S��*䧳5��:�:FZ�A#�:0�r�������c��@B�HD"���6E�W�Ew�!�^Yz��a@���=� -�>Հ��7n�閞,-vܣ4 ���D���|�����_�]�1?o'�rb)��fv�S���r5M��פ�f����61�UKF\��E )E��x�Bc�'$��+��١jaK���'De�p��%�F�l`x��yj��\nɬDK���E+pS��샦�?�8$��	��)����i��EQҚ�Ud�Md�i� �ap��>;�۰�:�Ǹ�P����!�)x���Af[����(�&E�����yJ�d�����w�^c�Yhyv�=�;$::5c!�d����ثR��尡em��!���K|1�9���у^���)-o:��&�n������H�)%�Sy'�ؔ4�*^n2i���#u��Ԁ͕#�p�ڂ+�$���-�u3r��^Se���Q>���(�����V�z�zK<y-h[���D��
&�r�qa�ڈc�$�fd�tKŏ�Jܠo.�`Or:L�5�Jv����r���Gcϟw~��S)J�#Q���
����:~G@*y�B�nP��u�P�,��t��q���ˇ�}=���G%@o�=���2��I���G��;��n ��h3|��z=�˲�ϊ�vF�����FY�O����kY��yB^�
kU�.�\�G���hi���W?ne��h�@j}j��i4����XZ�Uܟ�έ�E.Pk�|�g�����T���+[Q��+�����S�b'���g�D��(g�\x��9#��/,��!Y_.�#Ų'�wY�����Z{��d#K�F���ߎ��}7x<���� [l%�ٝq]л5����zfZ:����c.�p�p+�|.S� 2�5A�(\���$�vaf9|E���(��}���^r�1bf�GF�1'��&�����֮Dw�<���C'a4|o�oJOh��^ca�����1/Pyf66Ơϴ����%�8��y���f.�;�}y~��I쳼#M`��"?Kk�b�% ����Աn<���p墥��CG��L']��[ݬ���O�ec=���D�@�O�������k3���� �����/�j���m�����T>jc
3���݅s۩~I ��4�@�QF1ғ	/k�9�W�y뀷��1k�K��pY��;Y��t�P����P���Za�\�8�F+�mg���,��H�a�Б�˵�m�)s�5Y�6�.e���hu4�"�l����`|o9Gu�5�^���)\�����k��I'�	���B���yO��~<qIݯ�zge%���eU��
$P|!<fb�F>�D�� ��`����d��ҟ82f>�fR�$)��C�V�����G)��w@���?_n/�h��g:{!���5�����ZBlP��K@2�i�:�<*�{C_M��*TCyt�"�`�V
������<~�U
zA`W�~I������*��=�&��D�"���z�eo�WjL��XY�B�[�ڞ�m̪�^C�Ѭ��Lo�2\*��o�M�#�f�VZv�@7����V&�������́�~ӈ<�bG����>��gva�c2�E�;� ��$f�b��K�B�K���	r,]n��ޅ���XG�^���a�?�?8�Z�N�a%��j���];w
���q\�g��!����*�5�o��I��W��AG�$@��M_GR���y4[#���6*����og����9�[�%��qr�t �i1	ҙ�����`�9
��"dY�y����cfW��+PMmQ�P����`� ��-�Ұy����y�����u�;`��'���*��6⒟��oi�l��x#R��2D.j��x��Ͷ9����%n��8H���=�Xg6�x2�VV�Őy�H#��a�"ӿ�vT�0���(�>t�d���.,� �dl�P�ᄏ�����+[4��FQ���jPu�C��'�&�S��Z���Z�Ņ��1V-�/�>Q�^�*\M���˜��̠�����d-GA�j�.I��73��։�����ǥ��w6� v�
����։�5�8x 蚈�d����﯎����A�$&\䈐�y�x���M�<��?��E%����1$S�q�	Z�6!�s7��-���DO3���=Бx�ؗ����޺ʝw�ݸK�{�Ԩ0�D��x�S����Gý�r��$�1@��q<Q�����V���%�++0�ߴ��ꠈF�Z�;Y,#/��u��Ȏ$<�Wj�4�JL��Cp��,�\���O,*���3*l@�|��n_��׽З{���Պ�`gv7�)�a@� [#̹�V�����fg�N2�E�Y�W��Fr�%�>H�/�6�?b�J,�o_�26h���/��!C��<ͻ����+Q��G��Lh �G��O흨���s�H6���Db�|�t��8��t��c�2��"i*b��ޮ��h�P(S��J�#���W�+�-����B�?�\Q���%�4o���2̿?�Ւ#���:�nig��[�yd�4�-�D��zW��!�SXJ�o�� t�n-��Ϋ�$���pC3c��ݽ� S%���M�.�^�������� ��}��)Q)�jg26V~�SE�"h��6����X���%�����E��R:�Z_� ӎ��7w�a��`�]>�b��|���_-�����K�����xە�ǛF9�A��Qϴm*��<���sR_\�܇��\�	�Vh<���M�5�m�A�C+B��IWy�D����	��)D1>R�9)c���r�̽���p�@��s;�H��Xґ
�R��N¹�G���*yg��'ɘ�	�߭u~F��ވ�8ުl<�H�s��:�c���u��
�*B�bP��Ή6��3�X1�9�AIj�eQ���Z \��X9�x�1��?l!���	���g���2�1ŦmsQ�k5���z�I
-�i��l��koW:�]�b��c�i��� ���Op�4w�c���m��i�&�ME�b�0tAţ���[�&�q��;y?q�E�u�l;�m�������I6זo�pXR{i�J.ӸZ��p�_2u����38�g�\�Ar�;RW.�-֪����IQ.F)�����O��QN�d���p��daK���������ų{6>�nM��[�q�����X3�M0X�'�1�ſ�W�Ωנ4�[��7k�ڣe���[��w���u��Zؙ,#���C8���=��r��z��K%��ڰ�r��$ۅ��6!�E�����c�� ���j_=�,��Җ �1j�

-�edH��W�e�6C2 ��F��?��#��x�/B���#yc��&4�3u���_i~:�e��g-r�m]�|�M��b{By�D�)��b�M��Wrs|'!�3ƕ�l�B�'M��	5�RbZ~,�][��sm�ɸEB��rf�5��6�46�n"����S0�^t%��~���j/��,�:\~��	5Ap!o�T~ϟ,�N�5�`��hA��(P�|�b��PD�P��d��A%���>0�л� ə��O�5�{���'i�/Sr��	���唼��Z$���-�����yC�'I
��Dw�<)=:����ga��gEr�Ç͞�I36�b6��ڰP�
M�ğ[c�}�l3�Z�x���e��Pg�p)#������~�/���2�&l��R�qB]��-�b�6Y+Z������49|r|�D#�+Ge�7|����sw��ogr�P0��o�vu[��*����'�k1�����TX�| �4&b��C>{���PP�	q���ɦ^ɞ�^�uk;��S�=��nf0]]n���{-]�f�r�]4~x����w�	f����tvB���:��Q%��%,)�(zQ���hi�ћJ��ȯ�p# ��E�����![>}�� �� '�X�<���PUM�_��--۠5���Dˑ
D��Q*���[*�A��R+�����O����*��i�������waP�C�&�GkpK�9�0��X��#�iZXX�7�',��p�z����`��ø�f��n�|!H?����&j,*O?&���JWqsG�>�T�� �T3���1jC����񑴡��}�y���+l4cGn��=w�e�@�R#M�`O�����ל)}�3��9~�5]���ބă���%!�K3l�]������D [�3��kP��)�E�V짢�kUD��o^6Ur�Y�2΄I��3�R*pփ$�Yo�j��;���Wy?h�-3͕���}�#�ڨ�������X��2�Q%��V�.MY\��������C�npË�J���U���)N�r�K���h9iy�ä���P9%��d!��"1V}��nw%^W��� U�2���+>�s^Y7+"��Ry�U�{�S kl�MԠ�ګ�S���VK��baC#��e��Ce@�D����,ZU(�@r��H�_��T�<��+���XG�E� ]�o����J�
��\!ε���Sn��DWXQ�ۿ�|*+�d�咇�cW$�ϲ���vO�����>���o�_p��D�LT�N,�?�������3��r&��^Jb��?b ��źe$8�a$�hh����ޚ!�q<�K1^I�Ϟ�5�uT�]���K�U9��6w�׾�"h��K�X�֙CǼb��7���y9��dz��OK�фV+�>*5hz��CA�|2f�7�}�25\c���K�����Q��.{�CO�x�����S��#��r��p@��)��4�Y\���xsU�dQsY�$���mVqz������e����BP����"��y_����_�S9g������4�8nIF���Hs~V��
#�V����'nۿ'W�,uѢ�]ǁO��+�Bu�	��>�݅'ַ�qWØZ�}QQ8��,�l%9.h>w�hCNA���
�!�@�	�+k�l�(�<�{"���v����ԛM]J@��ŗ8:�	f��n�������C	n���7;"�'a�q�?����*��'[N�������r�b�d�,��*G,s�?SXFw�;��2M��S2ev[;H�<A�����F�^�&|C���)�r��[J+�X��_�,��E�me\Z�NȖ-�҂�hY	u���_Ί* �/Am���I�#SI�K/$�ʁj|�w@�g^���;�+�:?ه��@Z�L`���:��F�;1d�V�|�ì��(9}�Biq�>�ɻ�8:�����9�c۵� ����>���a��a[]���x]T�����yF-f�"�WX�o�����2��9@�"q(����C&[J��xP�T���L�6�����b�&a��>�=��.˷\*]޵w�F��`<7�G�F3Bz^�	/�	�>Ch�Tb�p�xp�R����u\�^X�&&P��լ�)�@a�ڹ��7�S$H�d�@m�{�[�p=Y���BⰈl�����CPL_���fXb͓9�\<��g?�8���N���'���V�w���O���"�v�؉�[�|�RRˀU�w��N����'O ld��nُ�|'?ܿR��������W��J�R�S�ӿ�n�}v�
o����<Q-�����v�\��boԞWu��v#���?�':��}��>I��^��r&�)G�����h}��:E�*�(�&��C��JYt�Vz�����%Y�hΜ�,����V2������
( "ɏ��6��Th�9�N�e!a�Z>٘�p�׹�	�^dݩo�B���.���w�GOi��-%�5���ja��Br��a<u|qV/ ��)W�J��}�#�����N'Lv���F�4�Y(j�u�5C��U��Wtcy�� P�?�Ϛ�R��Ν[M�d�m��M��PXQ;W1�'\�����c�0��WH��Z��"]LȰC�X�/i�Vp�S����8����@K��"k�f�w�O=3ߖ�dM�߇����qR�w�U��O�h�`1�� ��W�M~�*pO�E�Z�~�wP!ܽ�-�y�D�0��������&��t��Ӭ�'�p_8��@���)��0N�͖4�6㖃�A>ade.���~>��[ISH-��Ы�:{Ir�TJT��@q�#X�aFÔT�m)��>Y፞;��C�_8+`��+��,-�d�i�P(��y;�*��S �U!#s!�9gjS`"�B�7
J�O��:;a{��mJ~�E��4 dǺٻ�� F�������zQU|Q��.�lE�>w�1�ڟl�����Z%^ޱ�;1({Y%؅,@�Ҽ}C����.l��~�H�~§��2�%��pb�2;![ީA,")'i����2�Ԉ�G��2�!q�o��cOo�U�0W�Z�6���</��8����F�q*Io����.,i�ה<���N�W{����./�>�o*|4PI�M�-#�v��53m)��|�<^$�4���hj���SS�.�8���7��0R�T��*��#ەN"�-R�3Zy������
�y�w*��*�R�G���+I��c\EK����(GƛU�^��ևD&4�w�_g��pT���=(�s4Q�����!��an�r�Z�S/L=nB�[༤�.���k�O�%�7eZ�*,�`�ȷ��s�θ�>�Ռ����C&��Z4I�ˊD����z[�Jbݚ�Iy�j�c_L�̻p�>t�2fG�d��mX�f2�8� �_��/�ߢ�3�|:����%��+�,��/;�d�I+�.��b�ǵ����]$�����)c�Kk3�=���*-}�k�埣��.��:]�� �B�i�ib��M�N�X�����F���u���,��"�^��{���ő>�Qz�9M��������ji��^�k���Ui|1��g���%��"��(�M�Fݏ���9Y�sd����x`���z�U���]壠J��ye<�9��m7�k8�̊R��O�R���:H��	�/�6[rR��BӦ6�1�҃}b[g,n��<��Q4���/�t7��4'�H.G�n"��g��i�m�$#�D�<�Q}���u,(Q�i�6���i�M!����y&���<	����_�ٜ@ �-���]�m3;G��Y���r��?S�p!��7���""�)�I;�\�aX�%82.ᮔ�����o��6��BԊ������u��{��JHaں.⵪}�b��-�
gYRt�P�~�F��9 em����������ߣ�\(���"V�-vډ�?�i�*�C�X��@@�= ��{'�ӗ�E���B�J��;Xf#љ��
�D0�c'M�&����=��~�.����¢,�`f�ƃ��Fb�a@9't�)��*G�awS�e���;%�*�	D�% ���R��NHE�TyQeH�h��T.7���v!(0��Ӂ�TNS�TQ��\�1ҦSCMb8�'�l�r����=j���y��R2�M[%��#�,<�.7�LiUe�m�:҈�~z�z琀��2i��m���%t��>>�#��;pn�W��Q�U��#��$�[h<�Z��XT�;���%A����g԰B(%
U�6��.����"�$��60���W`���SD��K��,�����q��ۙ/�>Q{1����>�'Qy��QII���$�MO�r����T{�Y��Tv�
@
/[�i2�h	��C�Q&�"	�g��\� ,�"��������ۡI?���P�!�`,�o�'arxg���*����'?��U~�D�)�����B��l$���Z�Ĝ2o\�2eʾ�+�ݘzt���v_ 9ҋe�G2w�[q�'k9SD�c���VR{&$$�ژ6�!��	���YZ�\F����J���t�ڑ�,*��)<&`���D�d*{u��.�M9��cX����ء�D�pN�/V��l�/�5�l�]G����ݥ�e��ٛ7׸�
]\��}��s"]�����q8`�w5�l�=$����Z�U��j�G���3�]�q���)C���Nj	�˘�/���H��m�m�}�'���U�!Whw�r,9EI�$�� u����ۦl]��ݺ��y��!��%��~��w4x��VO��F7y\�n���NB��U�N�W\�&}�����Jr��(�ǧw)�,�^l"�cH�>�O�s����>�ӓr2H).��ĝ$�}�=�2F�%���_�~��H���]+ ���y�v��(�%�D8I���!��9��i4Ţ2��i�\f��DI�B�"�d��Y���a�&�ױ$N�aR�^����G��O�@�zD����0��:.�M$2T�҇	�K�LZ-����E.*w*��4sP"�^m$'2]�?ܠ��G1n5���������FWܸ���2:��[
Xl��@O�C�XE������\�d����?���Enյ�)
�pM�t�lSF~���=y��5:�ӄH㢚%x	%���c�� �87/��:��/&����M�w�56{E/��r����V�7�[(z�(���l��Mǵ��ɓj�?�-��+S'�3�_8*TVU/4H6����ҫ}��gan��lةDG�9���H#�óD[���,�_7�X�����Z�sθ3�*Xޒ˥��E�+2��/����˺�!���� �:c����V �9��Uk�B��zQ��.���VD5}��a�9='t�m�����ј��m[v�D^�y��G$�� ��\����Y�.��S�=�(y-��E��+xJ�$xee��%0^N�=V?���7�,�1��}�AI౾�ɏ��ۢ=��6��#��y>�\9{��z��F
��ڪfP����>�4x4�G��A"�Y��� ]��Ec��׫�=�#
K�Q�1�J+{J��w�FI�!MfZ���z�i�ѭҰ���y���D�W�G�[D9���M�h�N'�@R%����s��F��8_�F��:��Nq��Ps��ڈ	��Pl�K�������AZX2BGL>s�	*����SgM��	��<$�=S٬(��a�n�zhں��rPW�d"�'��������V��8{�U���˴V����Pq(�.�K?�stf�W�R�M[��D��_y�s�m������<"B�f|V��L��g;����9��>�Bl@~1K�� b��x5�{�fa�����!ߒ�"U��j1��j�E� �F�G���3���N߉�< 4ۺO�.
d��r��˴�,��0�ݵ�kq�Zg'$�T
N*ԍ��7��'�^=���Q����5%#�g���X��,�-R��JL[C}��79n+���,^Z�
01���ưnM�!|����]�PIIQ�Ak���R
4��4�5���$�Zr,eؐ��@`R ��6T��rn=5���9C�Ҁ�w��C��4�2��+������7O1�j��Y��a��E��p�x�|�
!i��!��P��D�����F��m��}�Q5~IY�7������3���x?��ޜ�������_Q���H=J��΃4�<���m����r��n,?�����`䯓�ϫ���Mf�#YT�?b�E���_�@�,n�$�=��i 
�ϻwp=D)�g�E"8���M�ǘ��������ng��n)|��Ump��r���K�X6�s�QE�5M�n�L	ID���<��3��z����%��՗҄=�D�<g�=h�����X��HJ%缩7���~?��30Dc�{aW<r[:����+�KZ�����V/���Z/������w��\%I/��0��]?���Q���Y���>6;&�/W�'�l=�79��
�zLvu��"?�h���މR,{����%`�ŔCwE�ԚXci��.��VƄ��Lɦ�NGxé$��Rzw��Q~��vW�<�CI��3� �m�2/@'�k�L<�o��9���S�+w"�-�^[���׫㐘�NĊ&�K(�t��5�ըan�޽vǓ���S8B��p�s�!������-(��������t�%A��s���Cf'Q��ף+�AX�1���=7��&Q�ЌAq�˞b��?	l��(mz�(��Ø��J����el����o�b��m�%����-[�{��[��8c������e�gbl�#B6*�H/u��#�Y��GRa��V!��SPSɦ*b��u}�&~{�2�&�-��._,Ar���	�.�ҽ�ɟ�s|VeɬG��u��i�/S�J�������;�@@4}c
S�ɴ�\C0������W��i��QQ�0���K �(^��A�XD뤎�ug��+���'�r����ID�mx�/����7�T<������0�o���C�/��k~�l:����Xe4�G��}�A���p��g�гΕf��G%b'f�VC9�(j���,wr��}&����,�sȎ�0�XS�P�ED$�+]���/�z��ngB���l~.K�A�ߤ4Ss�g��[�[�e5�)��O�@O�N �-�l�'�S��ϒ��@V�'�#�n�p�Yj5������U�~��T]*t1yCO���A�C9(d�hB��bP���0KG��"P�)P�/�]0���Lna���7Vʽ�^��6�/��|AS���}
U���3C�j�[D�S�i�Ħ���?��gR�����é���m����du����QފG�N] pf?�?*�i�Y�����1R�#��*�D��Z������)	u8nM�ğ��2�y��Ll���<�s5C��QK�z �b��=�ނ������z��+�e��0�.��#w�NQ/Y��t"�����[0��r�X����
�$xv�����}�^�6�è�Sů�O����Cʲ�3�W)�B��?
͚D�F�r�G�u�r�5�d⎋�N� �=�E�~��7�0lxS��d�(�09u��(��~�t=)��~U���v%y:�k)N����b!��%TJ벻z�8�]���k�|�[��69�R��E��5.%0��g��r�GR��U(���GL��
[��L��Ϩv�T�� �K�ʯ譾O�y#ʸa����7�ct��b5'�2N���N��yg�OK1�x +���jM�`��LY/z�3�u����<��d�w�[X%����6�����}��}Fl��Z��F��2Cf�BІ�.�+��>z�^�Ν�{y������`Q�'����9i2����He����O@�
E5~�/2&�(������]2��^c�/�dq��!��m�r�����>�.m-�P_�	gbg!�/<	Q������Ie��]`�Y�y��/f0˭<�	/KҸ����T3�)���]���<C�M��:'/���"3�n�A��B�tk��q�LK���$�����{l(���lki �I�QY��ъp�Aӎ�w\�"��s��j�_����8J}3���g������4T%g��J���k�KCy�8����I�D(�/.Y!����D5�N��{\�	њ~�%�GK���\`}V��Eǿ̿�8R�s�
�ױ���������o��^P��)\�I{(oin�����n��&p�rF�XN�(��Z�+�H9H bOݙ("���9��Up�# %3J�����&c�W�M�$.[��}a.�P��R�Ch�ƹ�q��c+��s�u�Q-w��E��	
%����jշ)�\&M����j�C{�b�V���.�5�n���y���$����f��{��ت�>�R��ǀ����KD���P3��?�4@7@q���Ez ���R㸧�Q�o��b��>j�XB�R����!qmL����◲�}
_���� j���tx�diS�\�0 �1���d�����i=|�"�G��������D���1��/�{�d>�@ȫ���-f��s0��;'C'3�Y�S�+���yaF�}�?�%Tn�'{���������Q���ݞ��>� T�N�����f�h��ěT$E�Wk	X�eD���Dr.�*�$�4K�����"C��a8~7�<]F��a�"[6��_�P-5=��`����iD�<=��i3l��Qe�xr��^��-��G��ٓ>?J��sGv�#��,\1�2�d����g�K
�2Y��ܾ�2�t=����W����5j���W��K;��P�hq=��-��pp�2�	�����[>�Ja�$0apL~W�Q9G�#�lF�e�R#�٥��C�3-�uf���?S���3bEl*y,}c�:��G�5���\HM�J1Q�t��J
1��+�:ǒ�mT21tV�
���O¡|Y&�0�9,S%�:�t����b'�(�����'�.EQD�1�����;�2�`��3� �)ߐ�q��G�*X�� w;/U��!�1�r���!���D���[ˢm�KŊ��,���{c��XHX�=d�zE�8�W�)�bv�v�Ջg��=QO��U`ݘ�*�
�]�E��6�I��i�Q��8,k �Z��,��	�L�Ւ���g7V��Fuy���:���U�����&����]�[$w0I��h��,���B(�l�f��E�P��꼥Yv��d����ꂅ4H8�YTP�k�",5lG�[�DqK��p2a�W	Q��B�GR���e��Sn����8$���ՒlacH��uElE�~-MM^I`e�=W�	&'�Ԓ�"��M��8� ���2G(#�F��ۤF�������K�Y�}�c�ӝF�h,�0�����%qf/�f��7	�c�Y~0��[������g*+��:�|A�3L񄉜��L��ƂM/�)����2�1���Z9���TG�|��u�)fM��Lu}���!̱���\F�8b����ݛ�rj1�I)���s>Ez��yC|+��p\�s���{*qH�����}F[1��}���2�l�=(�p,9�o@s�[��޼T�wQ��H�4�a��u_�"8ݯ'�������,��c��1^!�,������sl+ٵT�K�4�2&�*|��5�&h
�Ǯ���O��K��7�/2�}*Mv� �l�+DDA�0����}6�����cMB�l���G����<iݕ��?1�D�B0fJ����.wr�׼I��&ho1�85���F�k��^�}0�kP�2oQ :��Sf�aN�ne�3���e��i(�y��O�R�\{wЊ6`X����k+���:
:K@[C�Ŵ�A�Yj͒J�$����YT�@�>���T롖��v�*4�8U;�j��Ȍ9c�&���-���d7aD4L������J��B�Z:��t|!��=�#W�	��Ζ5#��j�V3��2[���;�=mgN���m
ۣ�7.�`�>�2��A'bz@�ko����g�~�����?�<c��+}��)��n�P<e��Q�:S�ZZөZ��%���5,���pџ���wr1>w��Ȱ�Ԅ���;KE�0�go���-G�/�"S��,6%��G��`��%Y����l�o��<��埏��/��3���,JA�h��O��KJE����7vo�=�����cF6*���e2��=r�C�Щ�[�P>�v�lŸ9�v�.*Az�K1���5>\2i\����\^1�V@ZU���RJn�����]	
��9�O�8kF$V����4�Ef�?����8�n��tUc����B�8u���J>���$=u5��Q�c
2��hu�ל;���lc�������eI�d��ri+f=�oH����s;�����4s�T�/����L����yy���w�.���I�s���L���_8..i��|˙;)���Z�H,�=a:���T�h�+�m&{�1��yhK�>>iV��<���(�{��k��z�@��i]�+c"�
�gs4��|�|�^J5��g��BF��?'t�PJG���,P_|Ȑ��j{2�R؛��I�e���%;Ԭ:�� (�5�g]�25 ����a� � Έs��)+��ͼve���ANm;�MQ��9�|��5�~�b�R�郶?%���Ќ�������&���;arv9vMv8�),m�����FwO�d4_���	�;�Ϡ��X��!dȲ6��{�������\��������3,)��dβ��Ʒ6_��9�uLޯ?��ÅE����.��e�\���i�ev��L�����#��h�'��9��-%J%78f8_�ˬC}SPƣS��P��H����m��V�
��R]Y���+�s�8��O2q����8�μ�ꮼ�]������7t-�F�g�����~+Vp�
�\��w���}N�l�ß�<���3��g_����9K\Ef)(]�E���GT�&I9 R6�I�,����!g�2<wl����ʺ?�>/�����8�!�ΰ�{pӰQ��fK/$c:YHRh �D��ߺz�'1k䤒dK�%�{��&��/*�$1��M�:��c��Y�Z�>-`-�>��R� �=�Vo"��jʥ�Pa}[�WgN�Q�iX}���Iļn�Z �g� ��/���R�ovy�U�O�o��s�DeT6�V��/��+U�����
4J\!���hdㆁ�_�Ĺ�5{f��� �]h��;CP�X/��'{u��5��O���NQђ���|��u"�o8����#�Q�ݰh!�|��qH{#	��vd�I���ˏ �] Yxk n��� �眄��e�����$�Txac�M9�l-�A����s�����MK�����.�ް�Em�+�%nV-��*4�f�a/�;v�\�vs�n�pqe��'����Ѕ��"��	bҦ�@�v�x�n`:R��r�hW�
�1#��G\	/�S�`�Z"��YP�?]荈�	�&�@{����4SR����2��گ�J9!�u�Q�lZ���%��F�\ᏸ�֩�o�r�p�`�z>ׯ��n/c²���ޔ�`U�����C��ID	l���cVOj6������1�N��WD���Zu.�Fx�4�G�|o����
�9�v��u�.F^��l�b�%��oeg���/~wf������Ѿ5���ƻɈ���H<t7�q�l��s�gdY�~���"�K
 �h����M��b/2)�̌-���A�������bL{Ap��$�x� @��С�;L��ņ�*V�gv^з�w-��V��U[�W[��P�A%�{,��<J��Ԋ�9a`�"3�2�{(X\�{d�̨oYi���3�N[J����L���)O���*~���qXU��ӉCt�5	y.~/���D-�by�c�W!x��V��\�c�6ɳ���P
��с�X�ߎ�2٨h	2���䈭�jl%<�pb���	| Qn�c�5J�/�}�=*\����t:%
q4�.|�?h����'��G&��~w0x��Զ���G��t_2L�1L��]�O|�Baj!A��{����u�'r����� �̂�E�ʈj�l��">Ϥ?B�DM.����A�v\{?#�]��o�zE��?�å/n
�g�@������K�91N,2���7����e�fB�2��+pn=y�I�,��'�{Z��s�Gؑ��>U�� 3X�Y5�}��$P�������\���m�C�i,6�n���ˎ�1�	��B���
]�N*JW܉�wUsy�lm��j'�3`sٙ2�~M�n�ey��a_���rm����z���W�j��B�u:*k��_]�<��r�����7R��|Sϯ�)���k��%����� �2$�S����+אn	@�L��H�֊��=�s��L��-l�r�b´<� ?��;��_9AH���3��iM;�;���14����*�50��9k!����쳏r΄�?z�uq�Z�1��n(�H(�h�t]�ح�O���S�t���G�oN�;�|�0 �nG�Xr�'z�,C���N/G�_�TI��e�V�=	�g�4����A�<�7^��"}�$�ED��������H�+y��L̃��&�ѕ����ٙ�8��z�lE����c#A�����1Nq�����	.��Qm?�T%Y�:Y( ��D*���� ���}�mv@��6x��r���4f���a�R��@GY@ N�-��n� �(?h�9]wcQW΂F�V�����
���T�3������k�F:^��|�J*L����F�z��{�X˄R��|��C���P��$8��|5�`���TA�Wc�L-�c��MAu�R� �QAA^�'�Iv�>�)�
��+�?O�qiV�� x+�:�*�Yd�b�>����V��� =�����)��7��;�ؔ�ϥ��L��J���$���O�o{��>��n=��>�y��#��8ei�M>�`i���H'�/�q
�V¼�� j�z�)�v��#k7Ǳ1�M�}~I%���2�_����Y��gL2�9Z4��Z��gr�Q�L{D0��B��|���̭0�B��+��I��'^���i�g�K�(�af��>D	s�jI���>c�/��?AV*%��8m^�]��'�6�x��\ ,B�]�'~?p`����M�xX'-=j��m|L��v>7�Bۜ�w0 ��y@x$92�)]�\֝saG���M�ƌ��][��#�ۈ�c�u�#ӞWK罓�ޱ+���{�P@��Q��N�|,��@(|vD���o$� ���d!�v��
�>y�)�ז��i$y�+����ԃ���r�E�%�O�叄�Qc壀������ ��1�F9�vf"���̒INRFMh�|��0����a�`�_
�+����ヶ9Z��0��>*ԓg��Ku�L}��q��n��o�i�V�U��p`�B�Ӂ�w����YQ�|��+�keBU�E�Z]۝Hj.��M�WC҆�M��v��d�-&'�C'����(�--�U��Ț/�_���+O�?<��i4��3���RP�;$�b�P��,#���v�\t��I���v�<�P���-��.�>Z���/�ā
� 2��=\4}�ȱȁ\�tȫ�D�p��3^q� �*���ɵ#gi��D��$�sj���A���ʃ�L��h�����d�B1Ao���R�b�����m �Ǫ`����B��a��My�����tvم��Zf����V�	��2�%�H�:͝N�̒ ����gwʷ[[�A�`��!�C �shk�����»-����2��>���U:���m��?�1V����^}�+�>�_�IE�@f�$!�}��ؒ5)��T?A��'�D*Eٝ�a�8��r��Ӫ�A,�1!YbTXU��,�Ҫ�vճiPR�3UV�^)3��k�	�57��h��3��̏f�x�>.�>M5��[�I��r��@ݤ� �	��j���g�f5�ڇ��B���@ua0E����ټ��D4�|K}�a�MU�G�=3��	��{��������P�ϴ!3%��-����)n�8H�we;*5�Hd8s�<'0���|�P�/ŖM�\�Qyq�:��Zs�,C-����0�O�\o�<0&JQ�h|���'�2?\��{�9���z=���G�rr�7~�2��7�e(D�CS)p��h~�Y�?�Z��R��v��Pi���Uz��k���8x�����!��.A��p,!	k���,�e���B�b����o�V����F�����t���Z�5�!n7�q
k�-��n57��*!zͥ���BS�5��&3��m�K@��\�U�㘁iU%�,�v�f���`���v��@��y
;0�,o�]~ǰ�WT��60r{�̈�x�8l@�
�����.>��O�W���C�y�_�cfBp�O�u?�_���|$�<�.LQf����E�:4���a�n\�Eq]a������'/�Z/��������p����|���wUƉ}r���\�=�,&z���w��z�#|�5�����\	)G���tAG~�PO�Ȍ���U��q���g�Yq�TE���_0m�"������'n�)��K��H�{�Vu��a�#R��.6��;��ĝu�6zR
(���WcG��ήDB�̀�_~@q�'l�Z1�7��"��r��RǱ�@H�6V�z������:p*h�;��ʄ���G���ǀ��W�
�G��d�(#j���i��M�DV}k���ۮ�G�Y�*C(ACA��yt;�P\iJ�P;��Ʊ��ɥ�I�)^�8�sm��	"I�ĻL�S�b��9�W/���]0��^t��(�h%�ru��r�r|*9��q9-bP��	��$ui!,��,��� ��pr�6�C�9cK��C���!g��K���5g"�O�|��Ғ�[�҆Hk�M{(M�`VYa�ߓ̣���j\�w%CY�3����~��ʫ\� ��W"�~I���w���W	��%x5���l�N�`�k&����viȀKr{��0�N��5vedGQX�%<��t��|+���L���AǼ�9���ʈ��gn��7��'���Sj�3�AZ� =ׂb,�
@��6ߪR�irO���S�jB�X��i��.kv�U�ә����P;xQV�6��J_픎�e��!�no�r�h�����N
�Y)U�T��Hy����UZ�F ��?ݻz~_�a靮vMO�]�#e��Jp�`��r�$-gH��\?XU�ȯ@b��8���JNb��c0矔��^��߇_b���Z3���~��b�"���X��#Z6è���5�}kD���_�Ǵ�`�>:�xXOA:u�S�N�,H�����|�=��q�<C`��P�Ѭ��]�<�{�R�CBR�0�Iwh;�X��1�/����c��1w��2N���)��y������ͭ�6S��A9]�L��r�������I�kQ���N� �����Q\�׻��?[��G����"�.Z-`]�0v�j�)��_]�
\����8��[XH|�r_���������2���JU�=F�kN��B�[���v�����8��^�Dr�P�ˁ�j���w���F�Z^�������6�%����k�(�}�|T�,x�ڤ�g�����Ae��~֝�"�C�1�\X����@�m��<sA�2��'iRTw��1F#n��;y���*ίdrLHY��O~�Ն���3�-۟{a����� �C�I�|Z �!�"o�K�LV���]k���vɯW57����][�|�_R��X+���mw��m���O���;�؇��k*V�=�.��d�b�]6�u�K�	؊�f��;���o@ܩ^o�#����s �5F����!-]���h���Y�d�+��j�A}#�[a� �xx �����'1�_��%T�=X��Ш$�SBh�ؿ�W��x�X���]���.�#��^`[���B�}g`�g,c�{�L�d��P�[�c]�� ��O����r�ʴGE������)���<��!	�ÍU���,���6P���bD��9�m5Ŷ�Ћ�;8.I
�������t�M艄�4�}ɼ)��H�9;v�sֵU�ɥ� )s�
B{J�ƾ�C#�{ŗM�̢ߠ�E1�8�P]��`�����s#�x�ǟ�c������]6���į#����8]<��+}�Y���}��;M\��"� ���5��S��@�Zn�E�e�!D�!���ʹ�ƙ����ڒ�Hh B8�@|��Ո�����ey�����/x�������"M�y���o˱V̀f,a��	(џK*���/�����q��v�E��v�<&���ҹ>A*B�:�j��]]�#�&wV���Z�8�^�0,�@��$M{�Y�܅���l�����j[�C�R�}2Yc�9�vėpYO�vj�5�sp���=�7�B�	U�A�s����R�+���v� �\����R��6��I�Y_��&�,TR�)!�DޭX� ���	t���_hWW�ΠH���&�N�$���]���Y3����
me��yGQ7� �cO��!������c�����A2l�Q+�|�����i��s�� M���i؁/�Q�ɱgcbMhMsPF`�ӹ�+�����¿9��o��FC��E�V����S��kMk6�Fx�:��S"��Vf߁���\��@�� !��ߐT�S�c�z<���br�-_]�y\�I*�,���{j��F�C5;e�v
���`��}�jЀÖ�@]��R\�� ��F.=�x�#}oҷ�>��)�P�< �E)��(����be�3�G�{���ܘ���߱8t:?è���}46,Պ=�t����p�>:�����G�eT4X�$m�7�|���a����,� �
=q��g`�sn�m�IL�m�_S ��0x�J��V��R];�0N����a=��7���Zl {*7�W�0�[.�#Ë����z����c���ўG62�G�n� ��JfEOe�.If��F>��v�[?x��ix!Q�6WWJ �#=���=��D�� ��=�*]�^oX ��6W/h���<<�YgjnΨFH\�d]	�FU�����Oi���Ff�3����5�d���8�B����t���ǧ�p��
.�v:�&G�d岱������@�堥�2�:�r}2�Y�閳Nx�ه����!u��H�����^�EuVV�^�}nh�g��W���0�#D�=KXt.�~����ʱ���Q`��3,nD�:b
+!����R�+e��W�.���է��rn^]��ߕ�_!8��"�~����&����f�<7ǔ���D�A�8/Yr�G�U�w���1��F����|�v�L�d�K!�<,eV���!���M��1�P�E��1+&�y�.*u�S�[��Qpx@9�V
FR�Ta�F=���8m*��-���i��Z�ݲ��?$�y$�
�t�r�eʍT唏�����1����1[.��l]�m�8��%��9�?3����G_4+�G�}��DV��M�c����70i�]��&#1�r��"��6���˖�XOT>�"�Ck�h(���)�֠�J:�7�ɀ!?���-��z����8JM�������H�9��	 ԝ���v���J�3kN�P���/��y0�M޲���0�vsxN��t��բ���T-G���(K�<D�����˦Ń��6I�cE�h�d|k^
!N�vi����W^{�pp������б�螤�t���ps���i��f����*��Ψ�͸<y�S
����eg�mU��EK1���ʏ�.-e�f&��X��8��
���E�7
�u�@D
�\0ғD��ʐ͊14��j��Q�E��.�\zl/~Ĩʫ�b 2�l���H�c4�uH�O� y@b"�"�Txf�zηx��IUN$��M$��:�&�^ӆ����JJ���k6���D~��f+�yX+xf�`$�x���/1Ғ��dĊp�fWؚaGn��ǵ�ȡ��Tc��}����)��w�E�V2����آ>iC��8)ր��ݴ������8y����>����bא��3����$
Hp��$ED��*>��]��Ҝ���y�d`�2\�#�)ԛ{ߍl�B��ɀ��JRK15rKy�x��h`m����,HJ�Z�a�$N6�_v�}���O,-�R�:;y��6%�5����W�Հ���_N����旎,���Qi�O�&c^�޳��&���3����1n�~k���3��ƛ$��Fy�tlä�z'�!O5oN����NZ[C���0<v�+�B���5��J՘�@�e��p�e�&��(��a�;R��,i�95'B��+L��	V�z�i�ہ�H5�/n)鱿R�;t[�����WC���Ik��]�*yD����d.�k �=�'��RZ]8@��ՋAUwդf������'����<U���R�_a)�TI�#��?������}�{-����G�;�^��=pw�vyb<2#V�a��NK�n�}������D(�r��Cb;�=�e9pk��'�3��Z�ф�Jc>ؕ�@՗���i�5jx2���j9�w	��� ��d���`Ƕ�"}�F�{��[�
��d�oEh���v��^�%�.��9D��\��S����ߒ�2��+��5SG�E���  m#�5���7��ޕ��w�g��\�e� �1tz����䑖]0y�t�W�uAC򛥤m#NWՃ�[W�1���|:�C;}Y�C�&���)�^:J���y!�i�����P��l��	�Œ���.qV�O��<�$!y�!'.`F�E�����t�xk_�E/�_�|v���&�ϓJ���� JVҺ�w@��<�l+��Z��Y�J�E1��x]��yv?�l�74�[�����>�r��W�ib]�D��?�v�懾�+c?���s��R�}��W�ug'�oI�$��'g�,�����fO�]m׷�����.�GҐ�O���[	^����!:���~��zm���,s�����+iR�o8}�?����{^�A���X�%�+��`m,#ƈ[�-)l�����=��b��{0G�q5�$.�]\�l�A��'�
�&�q	��S�e���w2�I�V��HD|д㖣T^��k_�r���6�U&'�ɬ�43$�[ˮ�O���]����K��/��-�kP"�����O#a�z������V�x�w�~����e=�(�Aaa��[�%�
�\��a�-wXP�Q�ji��(g��y����đk7����By:_�H�Ƈ��y�_1.�;�\�[�o:�K�g�\f/�\#�-`P)�_�>D�?�PN����=����=z.e��U٣G7,�Ωk�i� �#�x)o.h�7������/��4�A7*��ʋ	 �W��u�G n�b���h(ŋױ� /X����:iyHي[Z�w�JD��+�}�2�@�Z�,���o�/�)����{���:�$O�!�A�\m���`��Z"�l3�rZ�%�s/��F�t��?gZ|'ֈ	�a�p�{/���/�~��چ�mI�d��w��J�����~"�~[`�b���0��	��f��L�<��c�a����a[x	
3�&<��y�k�r<�xr���fk/���LJ	� 1�;�0k@L	�ϟ�ɞ9�Q�|���s$a�޿)񟐗�0�����lme,Z�	�Uw������#���CWJ��t4⬝^���9qH�����S�>�U���!I�	y�
RFYݎ�ֺ+ػ��̵��K�a��-�	��1�,0�;�<,�p��u6�Vn���UdK]%`Ԝ/�t�O?���$p����&�$�`y����
�săgc����8�q�������s�-��k*�VR{s�Ivsg�Gw�?���?6ױ�)g^g뗷��c��.�\��ȡ/�����'��_d1M��4�}=��uDn��n���$��@�u�޴ΡD��� k�Ԕ� �m���{�s��k�<#�Ft<m=v�֏�Y�3�M΅����ꈓU�:��A�502t��c(�d�m�B�;���~�S]ь��th��O���W��j�l������{�uv�����k�TGM�4`�x�@�*X�����8ιi��J����g6�h�lXN}��@��(�3Q[-8�&1d8�������b e(�?���t'%�B��\��@~WǻO\���/5:Z^Ҵ�8W����hWVj�&��%�銦�F}�#��϶����A{��|�ȢfrՄ08 �D	0{m{,G(��<Oy�GmR��D��	��%+�I�`�\<�1��ߨ
���H
'��Q8����p5�zj���!8<���!�p�-�ue_6�@��Y����o�\�ۮˇ'�%�����QzCRS֯�m�s����N/p5�m�E4�lH&����·Mr%1�"yo�8�١h!�_����a�����mc2�'�`��g���%��f���h�x�5y��T�������8D����읓���`��X��T'h$���7OA���Q���82��#̈́FU��\"���c�މ/=�m�v��eF�h��2*�uT� v�C�C��?B�Ez� !�j���f������)�zKe�~�+ǌ������	�6f�e(:�� �;����N�&]��$`=VC�K�q(\�w� ����h�TW����z9�5�r�U���g�S���r�z��0�X�k��!�.@�٬W˪7a�Ԣ�$�կp���N��v�=��]�g�k�x�M��F��5�-/���� �0���0Ii-�]{mt�\��7�﬋���9� �в���4��Is+�Ȕ�I�wZ�^ɉ~�ܒ��|֧"�P󊠂+�(y����w���N�k5��`0(gc#Ě�����E���%N�3��%'W�����ܷi#U��S����ﰽgbj��I��A��eƘ�l9Ъ��Eݘ`���A�O5t�ٽ;A���[�y�"��C����H��@m��h�/��b��F �W�
Ex�L��2�s���]�Y3(���a��~Ι��T��i���V���Ϛ�o��1��ߑ'��M\�T��kL�i�	X�4j
�f��W5�IN�Yztl��� s�����w�ةg�<f�7��j��{O��h�R�Ӯ~G~�<��K��aL�z�J[�J5$G�����9�K��d,w��wurXG��ϻ4��Q��]U�.'v(���;44�F�Y�J
�����A-�	�L ���Ja*��}��g��X�_��W�>OիD��#V��W��3���M�RE�ғ{�X �NpC)'��Q�V�S̣Թ��gы� �NP�B������:���_�-tӆ�� ��X8���4B�xoV�$Ւs���;_ߝ�+��	"�?���j8X^,�U^0"�iŁ(�w񖼌�`��k��ʪ"N�$�/�u� n�"����%��\��~��4#��g���C:�H�<k�Axxp�ƒ`h�b�@�+�m�(MA�VK"VM�������܌�ZI��\�R������r֢�1/�:SAYq�_��]�.W��k�":��8����S�A���^�"Z�:�G�o.$�Y;m���+�� U��:#�7G��ޯv��%�����3�a]s\	W��b;��H'�u.x�A=�\_o�muʍSt��(�UT�Y��?�P����j.��e;�)FX�TQ��rQ&g�8�#���]T^)�,�ᜄ�1d�'���B����#'i)T�}���lu&"�|��dځh��1��%�rG'���?�����g�Ev���k"A3\�mO�M,�
ԃn�Ȝ0ux`�z����M�9�*eќh�$"IdF��bLJҤ�ZBհ���d]6���T���pCc!�	;]� ֪Y��GV���H�0�v�g�K��llo�2bd��{{����hE�zG.���F��;�%޶,wm��w���u�om��1�
����o�񤻚�_VdW��s�t!-x��I�"�-���FDve�|�:�S����N�8���$�+��~�9�+$�bA��[���ԑ���o��Z/U�q���>ND���ɟ��˕���Uob
o����c�{�o.��ٳO�Vo�[�c/��ܙ�����Y
�p����5��L��䍆��+}v�SjR���J�DB0n�z��> �؀��W��lRb����H>)��}�vH��~�Ql�V-R���u!�h�W�Ä9�A+�9W[�P�3Ęd��s'��Jme���'=)�� ��Uڐ���[<b���Pr�&��y6�2�*��n�iq���  >��T�V�U�A�?������ԥ݀��T��l� <�r0b��y�؏�P���b�6�.=�R!�%>� �>����
�&��?�~�и�<�nv���Ue-�+�'s��V5��oM��,�)(;�>��x�t���L ���q�X��Ak>��fTkk��s�xRË�#��H�<�󍠳����S����,]�	_��Ӭ{͠�M���:-z����i���芅 �l�^B�!�K�.,-X>�P㙻&��1k�/W��z�bz��V2��������k$�uu�9ϱ�b"��~�_t2jG~4n����bW&?�DP��'��c�:a��oÆ�oꦽ�>]��
��Q��A��]o���H���o�G�@(�di��(Cpv�\�����2Bf�C��&�B�,q���X�j�� ���2���ʼ]�i'���q��/�h�Ϻ^�Dlx% �ӭ^�>���!T��9��V�BB�H��%Iz!��# ����.^���}:ɭ�W��IcK���(��^t[.�W�w�I-=�����W�D�at_�����b����|��2�
�u�lG�V-�Q���Խ�z7(
M�����ߣ��,?�j��-�a�"ͥ�L�G��{_���u�b,�	���n4�v�m����␬�	�w�	��ew�*K����Ta��ۃL\����:\����;��Z�S/�Kks��}�� ����B�T>8�ɻ��a���������1� ?����ԼV:��*��F�����T"��'G�q���lE��`����"��؎�S".T����D0
�	c�ѱ8V����l9�Q��a`&���4|Zwb5�J93C���Oq:h��ֶ���/E48� ��9;���'���뀧�AO]��<�J�����3�& $�u��!2]O%����r�K¯t��?�_=h
,P#�5H��H�ظ�i�?L��3zݴ���M�3f#o'��aD�}��٢��x�v�e盙.�S%��0cw;Id����z�k��d�~��:�8���[,+Ҏ�3�� �1O_?��/�fc��pi���b�.��R�HÆ�ɸ�5\��7R���k�+T0ꖷ�����X��z*���Ql2�Y�8ݬ!��;ɹ����P��;��BW�Nn�=��\z�����Ofse5W��ל-�г\>f��=����\�2-�!y���7V|P�XQ0i|1������D�&,+{���G��6�1������b%��Y��2��Iޣr�/ ,F��Rd �r{[K��{B�ͺ�J/gK�?ɳo��C��`�z���Y���������f��ڂ��O��LZ%�6���������	�ɪ��F7
NV���JKk��5*B'�Eق��W�`�jvf���� >�����cBD�[[0Hʓ(�ق%��O�kۚ)Ȅ�����I�@�ş�K����\��iZ^3���<�������c�g��"~�`����T��i	q�ȅX�fMWf����L�'O�q�-,�3^)ߣ�4h�������9x¤zY&�]���;-k��e�ħ��X�����Y�_�+�������8��ﺗ����`�5������ 组��ieU�s'����D8�$�CT�8��.g��r��Z~�&����ÁN�Z�RB�Q����dT��b�b^(ވ�hL����6�B�ٶ��D��g����d*s���#qR��@�2>�5.���U���77~��3C�=��!�����n� 0HQ�B]���:gJP��m�W|�{��T& \91���e�M%����yQ>�������1n�P�Z����=?�XT7r� # �*���V9d@Je
K�ܧ
L�bw��^s�tc|�r�ϫE���l5)��zy�oc�!�y@�9%ǀ*��tAL��eM`�d�9�.��#qtӹ(l�5�f. ;�-x���9HO6D+oNþ�X����E�Ê�wpϢ:�npYL	����@�U��Fb7rU_�Ĕ�6�X٠t���K�.nw�d�2���՞��% �&�!x���)�L^=������G��.L3�~E�OX�1����*�gU΍�J�L�k�K)s��C��b�A�x�eيMvk��=2��a�:�.�>�� �C��MS�/]9��(���UP�ȋ�`vK/*%p�`ͥI^�ۋ�dx(k�
��y�K���\1�;m��Xj���m��e�V�c�"n�D��m��0��mW��c��" #���º�dՌ?�o:�#	��v��|��i�汅ٹu�d�-���9��hv��}�SZ�D8!꺈��ȉH���5��^8.�r֒��~��♖aD�pe2���ӥ�#��s=B|���cp� �s��^<�s���g�Je��N�@���6�U0SX���m���g���Kե�u9`��Ͻm�I<�.,,�q$�g�s�j�j�Q��Xӱ)�3F��N������R�s�}���Y/�T�e?��UJP&����Sg��q���WRx0'Y���F���>:)t�w�6K�.���m�]2zb�dE�乮/�6�;K.T�lX�Р$�8@9��_aHOզ���T����㺕� �;�\�JW=�8��Ćk?����W����f�f6�-'���C�̟z��թ>���z���C{�_ꩭKh90�e��8�y��5�)�A٫p
|C63#kDK��	��U�o����y������P˵��b��(�E�_��.P{�UزE����g�f�k��X/Ŷޥ��"i�͍��3���9-��r��>�?�g	��S��:w��h������r�XP�^�cH-�K\�!����o��3@{#��Mڒ~�}�)��y���R�9���!��A;�^֐��W��E��ґ���9�����S��[-�cL�7֦�RLѧ"n~`�P���RU�o��*�癨��sگab{�'Ij��8���	�j�|O#w��'�;���@g��=c�r0��A�����>3���0%jg�u�q) ����+��tl��zԭi�ۧ	J��H��)�c�\�%+d��3�ߵ&t�a
ݮ������-��b)Yޙ\�ߠ�S�p0�!"�&ʋ�eѭ'w"��0>4K���6R�w*y?�C�U�Vdý���h3�7b3�\��[YE�$FG�F�	|F�vp �k냌%����9�Ll����y�Z1��z�]�����_�N��w��d[�a.̼[�f��R�<��j�^����g�Y�:"�X������c0�
�A�J�DL<+ǩ&X��-b:����@�;����.u��X�~����N�f�1��^80w�]H�S��M
�&�E�x6����D
R�ӥR��@<8\db�,�%��=ͨd4��6�N����v���i�q=Y��E"� 4b# iTS.t�����@ ���R�b�Ѕ/$ED��~�X:n�H��o����K�	 �m-Lv�@��*7O@�� ��8o�=�?�3�P���������W��u��\�E��S&��B�'��+��HͲu0W�zJM\�^p�%f5� 2���[j��BɊ����FF�����d�7����x^eFq��e��j��ځRo9O���,���^Uc���ل2�&��ٕ?3��tvc�[�ů���%~��ƙ��)��F�J�ܔ�=�З��;���x��x����`��'����c��膶��L�P:[�N�; �If\AƍNp�Id:����L��Q_9A �ˣ?yUS��U�kߛ�|1c����4���G�EX�r)��A3��OtU����m&G!H��7,b��M�����[�ح{ V�7-�9d��]I�:�Aem�v�'��h��]��0Zc

'7A�_�>EJ�0]�)@���t����g�WE�!tM�X��"��E�6����BgSs�I\VŨ�x����f�dn�jh�8	Y�|�*�ȸ�7�^���'Xr�D�T�d�r��"���%J_�n�38ȴ4���H��2�x�qa-�'��|���Xa��ƍ�:Uq�#$��,�(�K1BޅwR��9����-�K,T���?�/p�F�mHX��uֻG�=���0 Y����T��>����ukq�ړa�=|5�$��N֨]�ee��GEYm��ኜ)|�9?!c6@"b��f���2���q��NTV�Yz�C��K ��HĮ�8��SC�Qʦ�O�)����CR�F��=#!$7�T�`�4�&��P�P]���aB���>�z���G����� ��Ŧ果gҘ3�P�%������{�5[2�z�|4�}�4wq�>��s 
4�T�?R(�y l�m���F�:��El�k�U�m�^���%���&rR�������}��A	a]a=�_�$�6���[���6:��K
�5���afM�|���A���q�Z05�4Swk� �i�z����%�W��<"3�yQ-��Q|�Ep���>��@�:r���D-��2��� q�P�
������F���Y�kz:sw�n��Mm��X���.��d5zQ#h~�NW7��V�e������G#@�Q�<�f�l��D�H�p1����?,S��&S��-9�=m��'��l���iƥ�S-fl?7:�>��̰��͍�v����1��Jz]�ԯ2=ؼl�!����`�QFu2�bzR����D�10�sk�{6����.�}�#�/\�%�*/4��2:p�n���p��02����jQ0$�� 9Q�!ap`���m�(��u��=+]�1�qc�]�;ۈ�C��ݚ���P�F�V-��iJ�QB�ee�"�7��2����| ��.VPf��O����	1�����	��%��B dwn�4����yGj�N�����c-X���}�_M�Ϻ����m$P��g���;�@ѝ����/���Z�4+�{�N�h,"��+H�ݤY����=�u��V���PeMS�Ug
��s�m�o~eQ�eRY������D�3�rT<b����3�Y������&��85j����=!�N Y�"0��+euMkɐ���L���IݻDE��D��0m�U�]K:��P���XLӄ�n�%󙹞݈����>���"����Æ��Un�y��rtE��q���<�ɚW���TN��A�8��/߉�\�n�T�"�.]Pk�0>�=.9�X�I���� ��	��T��~�>O�M�V �MU�ǳm{��bbЇ�sib���������P`�"X�I9�8���$�0{V�ڷ)ը|�0��Ltߏ���0��:�2}�����g��R���2s)��*��V8I����uj�QU���]��h�ݾ_��V�`ճ���a����> aa���7���	VyQT�y�gC����u5r�@޹��ԏ�#��f:��Z)B$��W@|FM�)L�Vk������?���Ř
y^	��}ωǗ�#��7ޖ�\`��2�v�)�h�%�U� �-�t�'�⨫�����	{�)��[�uL��q)����>�#y��v���O}��"'�\m�eE&9SԠ+�9�њ����7��7�΄0� �F(��kaa�\~�K�Q.Qpȇ��J�z0��5�#��e����񒹫QÖ��FoCt��
��-��|m�/����"k�ڀ:���Hhr�%��4:����
�+ ��=v��-���%_;t�������>H����q�j��� �}��U�����t(���7p;�P����k!�b���ֵ�H`��"��@1�
1�uծ�W2��v����8C	��5�G�)�*r$���9�'���f�8��{.��t�� %�1���l��$Ɠ�v���"����S��uҋcm������g�hi����7U�+D���Y�@�ҩa�f~z@!{q��|!�L��n7;.�-�\��ѫ�Wn	硾 �\=5UR�T�PH:η���GL����<R��je��$�`�Ř��a��X:&��D���d	j���݈��f�[@�	f)N�~=&k�t��Kֳ,�}a���F����D�{�����ַ��
�S�Az��[��)���z]Lx�����ɔO�5z����d]��@VH��7�pل,���&�;��K$�����1�㯜�ҧ[��(�3F�l��Q�͜�1pE�������M=2�ľ�j=�H	&j��g�����&��S��VKS�#�	*�ˋNu�l����Q�������8b�� ]=����S���ؼ���M�-���K$�t����3]SEp����E� s#�N�/�*��7�੎Jc*؍��Kt����@�GH|]���-æ�w�w��A���G鹍{=A������3�}@ {��jNe��+��n5��p4{>�����ob�>i@���3�q/���O&�}M�zm]��G�b.����/}�s�	z���+P�,��J�OX��f���I����Cm���5�t�c"��q���>��E� �,Jdw����Ƥ6b3O��K)"W>�lU��;l!���N�����%iَ�G.�E�f�m9���^���Cz��a_��]8�f~�ё����n^�{�U{����[u���aM}���9�+[q '�.O�ܐ�����]7ƚIK!�����P����F�t����~�W�^p�d񡚓��ɕ?��/l�<��`	Ro�;�rC���^u��~s"�gN3�+Bh^��W��<��e�nF�1��h�7�|}�R�[������	Og1��o�2Z^�b\�&�`0&�![�~��S�������ê�!�_`O>�X{p�-���D9�c�vƍ!�14���z������$]wD�Վ�����)�b&'c4���he�R,�j��ŝ�T���"�_�_[!���D^�$t��B��/��į���K���p��#�͂�� ��:���g��d���,+���r��>��ȑO֜�=��Ր�ĝtyr5���������6�?7N��}�T��i��%�g��s���>��V"/��B��q���X����ǜ���u��Q���>o&?�w�\lݓs�r�f�Xў��}B;Qf� ����������a�Sa�DY&V��u�Rs�ܸ�� ���Y�N�� 6'h>F	����Bh�u?�u����}���񐑪~�+���4��w����:��<_�Gt����Q��\����֍�qh;�Z�g��t�Y�0��r�[$6V>��LzdAT �Z��d̯΢w x�8����ȖY��|u��(q��_�	��%��Q�.`+��k��٨˭mt�P��"^�ً�����"�C��7��k��9,6�2�F���h��������?��o���q���\v�t�����ț�c��2_K�B�����?���*g�4T!�����P��ĸ���!]Gu*,_$P8W��i,sp-[��u�ɧ�z�d�W��	E�wo���<�� ��ԂZg��,�D�C?]y��ꯖ�� e��
��i֬�5[mh��Q��إw� �c��pA�)��:i���JQ8/S�n��ڄ���/��������kAzO,�Ұ�Z��s6(O����
��J�Yj���f��ik��9����[��(�S6ɀ$�}lh��55V\��������I���_nL#}�	��ND^�	��a,�D�Y�������-���s�9+�7�2�+�N��*��62��!@�g���"D�U��7ĺ[W��)���'IŲD'�]@�䚙�*F��	�4������ʽJqQ,È j��F�K�3�5�:ȇ.oj����'c	��Wzq�P���^!�ۜ7}��
4�g˺Ѥ7�eM�	�m�s{9�#c��@:�t���s��g����.�*-p����� ��.���S���n��J�C�Vw�N mS�%ڿ-)y���k���">���Lm�'$�aDw���N)�=��Q���hȁ��~ʆ1Ɛ{l;�CH����P����y�<��@]:��3�57�W���`H3�+衅�F�x�$JںAuLq�"� ���9�BA:���s�,/�ӫ�O�+��h�b"��"_a�'Wd��$c#�۰ς�.Nϔ�CG5����$U�@�l��р�%��a����I���@���>`�B�� �0 �	ۿ��׉�v��1�W���j���	��c����Q�$|5e���M;-��ݨ�	��(�_Й��5'�����S�/"�`;���:(0q	g���_Uݰ+�F�`�G*d4�u�+�Է5򱔴K�l�ȸ!�����zpܼn��|䓎	��/WS)�t�Yr�.��T����|�)��K�{:�����]�k�/�����{_�[E1�4W��"���� �A�D��r[��Z�C�ē�ʀ���<�	�,��K5�+�%늧e2wJ .Nʋ�fF��RXX�"u= ��sL<MP��U�7M��I�'���|W�6�X�mckP�B1�y>��-��;�A�o���Z��b��(|����XR���sl�BW�u�&���4a�ē>{�c�gb����ht,V"|���m9ǘ�ݛo���6���f��O���D�*=1���]����}��㸇��/�c�n֫n����M�6�$*�������Iu��k�i�b��Q
U�nn��A�\n���^Gs�� K?%�v�R��73HA�<�z�NG������Ɉӵe�$'��l1�d"�G�0+�:��/��r�߭���Y�$KhD����*�D*t���Ё&�6SI�H:��L��WN$*n�V���I�.C����qv�P0�`9�=fKĿ��O<�/أ�,[pKoؤ�Tr�EN�NV�D+��?��#EMS�i>k�m^�C3x*jR�e�-t|���=��`��~3��~�d��ѡ���+�-�}E�Y\J��]�Hq�#����WK[�]HL��qN��ޫ(�/s����$z��DŌ6nC'��Ъs��e6���؇U�U��-uaxG�TK�DR��(#��7�~���VyԏcJ.64����T>������%]W��I�w���&�^�Ѵ��ɻ>��kYɲw�4��L��`Q�lݓ�V��<�帢��.I�;صF&�5ae�{c���]�E��?�$��I�Ղ��̡Q�g��/8�`���|�)�w�5u[j�x&�ӹLG���$`�Գmr�y��8I^�1k.���87E�ri�G0�-7h����&C�0��6X���	����*=>��B�	�!�r�K�lo	{J�,~{R��>����ڪ(9���U@l�꘷+"(�r������:��=9H$Cm�P�=惾EB�%�qT�J�i0qI�N\=���GAr��vq����b�����&�I��<�濤��k�k(��E_�pw���c��w���+�cZ�V���D�-������Pm��X��2pP�
�5Xt��Ҙ�!�+��p{�^��]Ǡ��՟Cb����Cݧ	4
�,�8���� &a�";ъ�����)�]j��E�f�����s3b��U#?�8�9b�B���Oæ�h�(g�ңŰp}�k�o�&3΁�ؼ�w�_��>�s��T�:�a���A��1׉���ޗg��_����f�Բ�s~���!d����eY��:�jd+��j�����GRa_Ӯ��Ʈsݥ��B@��W�6�u�HML)/�7�ȉ�[��?%s%��/C�k��v��J��迢�
��8�<��K�4l͏�y̓�-��G*Թf��ֱ>)Dl��"gļ=�s�됚��mE2w�Vp��Ӵ�vS�-A,cD�e9��R��gg&	����w���kp����S���m��d9>g�����$wt�sw{��1!4��d�!�V2��P'�^ct�	A��[I�����-��r��?���J��m�<�@�3�@�Ǧ��s��?��q�0�W�j;�e5�O0g<���9>o�`�9��b{�uQ�R��wᷦ9!(��#��T� P���u�8��:'�R�+:����j�s��,~f��=Z�/l���誁!?�]5�����%si��˞׏1��ի
���w1�G|��Լ�3
!�>7��q�c湜cpVR��bY1
��8���q��pˋ(\�k��ZD�%�sI�p�Sak��5�!(��fY~���ŵ�?U�h|Q�u�Е�et�q
�5^f^m;���G?�c��4�ZrP����.�hK���f���r�F<�*v}�1ݙЌ[�iZ����3�_]P�"M�(���1�K�^���t����m��n��4�l]��L�g�6$~!7��# �k=J(�׏TO �Ϛqk�W�Mz
�W�*[����RU+lҫ ���.qons���ٵ}�2�H� j�i#g�����`��y�\�9p�+U���Dm+@��ͭ�S�����BUy(���Jmq��ƿK���P0&&EsQ�N���q�z1�xp�R�vV�\3#Gl��a̭3\xG�kKG�0�U��ړUc��z�;�j�2�1}H1%�"�&�e�	��r�R�F����e�(��Gr�PX�y�[��R�ν
����2��N��\ %���t����ג~�;��/9Õ:�㒤$��g���������_��֨�X�6{�<��Q~4�m��$ � I���z�V����MCێIx)�Wׁ��@���3�e�Y{+/6d����m}G�����q�"4{)�7��q��r��PR���&� ��o�����m[E��f�3���yyn�5�Ię��5�>�m�p��%�Z��-���gU	�����Mp��mU�\%��rK��˥��'Z+��[L|�FK�mVT�o��fy.�O8o�ށ\���l�7�q��h
�'1k�	E�|A���N�ca�%�>e�s
��Ģ�)�$k	�+�X�<~c���ǘ��n*y�Df~��%�P�䟱�!�"�Z�(���!�����z�FI����®oز���IB9i��\_+
�&�����̂r�8��{4�b���eu;����;܄�4���py�P�� p�
��*ѥ]�2��m�w=��=���<����$z�@�V<�h��oS_�$�v���R�|ȵY|+/�m�V*WĮ�+P@"�H���G�(Z䳠���j���kU<����[&O�[���	}��{1j�l'�ԡV����T��%hf��^�}!|k��C�+���P�x���O�>q{�%����߅���L��0:i�FbN�����e�lǢmꔆ|3T��`U.�o���bY�	X*N+��n���jC����j�����D��,���rHO�&�ǎ�59��� 4M0��T�es<(e�RYB��y�%��&��!Ok}�1���T����g�A�b��%E2T�q�^�W�!��1�Co�}s5~!咿=֔�>�-�<���<��wC�ڎa��\z(���֓�ơ����ٻ����L��
����|�}�@�-��tf������|��j:\���3�vbC.D�2�ȵ���^`�,�*޷ޥ6=-d��T�nR;���|��>`a��T?̬�0º��U,[� �\����`���4/3r	Q���wTBU�pxO%��ը���R�������3�a��B�QxJ���KyĞ#�)�X��{��DP�{���o����Ĵ��麪�4J�P�2_Z�� ��	�#�00���D^��ҟ���?M�vL�VN�Xӑ�xz��/�N5n�l�5��*zs� Fxh󳉓,zdH��3����	�bIo@ExZ(�����̽S69͞�I�CPb�_��)�c�ȡ��D_�cQ2.+�tV�YKh|�x��F�X� �37Oӣ�̤?�M�ע1L�}�A�n`��QD�7����ӊb�~nu*�خ8�"_�^q�N�߇�70��!bCt�J�CRZ�z�Z&%��9�a�g-v�_6�H@��1��j��i�����z�J@A�h�YF��Fm���]�~~r�M��
���+�b����E�j�~��O݈���$5oLe�a'�q��qq���u.����wC�����aN�6�����㴟nD�ǈ�<ۮ�c7���!�>�Iia�r�I Ko�\�G_���q��/Q:���v�q�!�z�/oz2��)��AWP8�)�Jc$Y_����	��W�J�%����v��<��R"8m��)��0`@���B��D#Π���;�褳������̹�3|�`�8��%�I����5_r�I0���&� �����{�����QGӢ�9eC��qLH�ז�=��O��a�NR7�O(t���K���OS���D���j�K`���-��f��Qq\JQ��мi1A�9���x;�pjm#
��f�!W^uL!P�&k��*02!	��L��O¼ަ�Zw�\�
�l��C�lgq��w�	�K]R�\�=E �t_��bC*��l~���}����\��"�Q��"z��Ax�r�������K����K),�l��S?��ˠ��~�؏���@�����*<I�j�IZ.���ٲ4��~!͗D��T5�W���=�i������k�9A�>��V�;_�`>Å�n������&szG�cz͍�?E��湅q��&t�F"�QWY=mv`f#�fZ"��������\Ff_�zvM�@�F�iM�Ć����ؚ)�y8�}�ْ�ۋ�
���u��F �D�K�%c��}A�I�_�d��ujN22ޜ���n�1pT�|���ǋ$S���� �u�%\ s�Φf�`�;f�](�Nݻr��R�
aֲ�o�zw!�/��0,��Ҡ�'
~�OG��������-c�@/�?ろ�:"�x3=Q�.�]�B�?�`���k��""T�۴� J�����ٻ:)BT�ج�<
���"�^�k+������RA�g�̣�����*���|q�W��+�H��a#��z�aņ6�iO*�-PB�i�^(�Ҧ��T�t+����u-����`�2e?�d}:��U����C��(P&Ȗ�H��,�p����s���O�~$6�r�uL�N��/��v=f�6�����'�"5�$k��@T�D�`�Pv!�9�!�,-���Px6����%lQ���9����h;ʃ^N.jӨx4�Ӌ	������v�#2�w�r�T�F�`}�'�4�T�%�T�H�H�K��6�>�
ޠN��e�[����ww��:���#���fP����+����m.�f��6�^�"Gvy��v	���NH\�̗(/��}��z��J�bJ�D��`�%��J���a����0��m(��#1�keG��A6���9&;�A�y�͝M�T2��y_.��gӜ���Ӎ�o�����=�l,Y_ϒ[�̲3[�i����r�r]����:~�������6PE�7Y����Ƚa&Î�����|~�Y�)����Jh��� }�@bQ��x�S���
�n,�_�֗���	�ڇNtb�E�9H[
�g���O��ْ��!�g�z}M�+�۟�E�f��0�*��}XNՂ�k�$J7H�)�8��<�V(g��l����6��Ϋ�(�Fy@2��As�<�Ȣ�	��q�Fx����!�_w���mEZRz��q`A���^u�0���P�jV�`{P��y^��l�f��,�V@���X�� Crc������-�D��[��(BU����'����=��b���TNH�BQ���k�t��41���0�(�5�q�-j�Ny��*�ZeccU9�M�5�g�ն�,��Iv��9�!���\L؉z��	��8��弊�	Ӟ�|�y�.��]g�H:���FNH��[�|:�X�	�s����Ͱ🷞dn������>���%��Yo�,���Zt�0�i�������b�VU��m=^(m��O8��Q7�M'��?u�Y�̽�>T�e�#$�����֯,���F�[����/����PO6:�9��R�喳�{1��������N׹���|���%pc2�y��u���2)�Q�M���$�E���������<E���o��j�p<g�kWI�B����o�b�*QtR���/���V�����^�Z��bs���>���TlÙ��}h���8��mj���>�\�~�O(z��(H��z.�:~���i! ���x���Ԕo��#%{��c��h~Lx����U:�7//	�\! � ���Q!�1�Q�kֳ�
��I����J�4y�S�?����h�XBo�N3E
��^c�q�Y[��	����[J�(�{^����I)
�������'�ɐ��j[����Ȇ���Bo�(�V�2_�����Z�q�.������7ZK��e!�[� u	��c�tIq��6}�f���ûє��P��w���^��L�Sz�A�2�͘����0(`���qb�gl(R�n�|���<��՛�l�6
R4 ~t�Y;ML4:	�Oa�)�l���	I��ک��N��a��dvv�%� ��U��$��Y"���h�E� N�ji�}�](���B���m�
L�����:�!�%����'�)鐳@�-Q?��u+/LqF??�h��I!#�/�q��E���5��t����IZ�:ZA�(~[/���ʗz�ܿ�P���+����[9֠���3iX:��>,B��p���xn��_�ߟE^&Jƣ\����=u��u+"���0�`{�}zUE��\���҃o�o��_HY�; ��V���9�䝚m�x��.'t��ŏ�׌�fK�F}/�w�\�z��2uz����`ȑcȫ)��x[I~�l�ca�9��7�h9CW^n>I[28�"ӧ�@��X{�
{\:��֠/;^�n��</�qV�Ŧ�]�擤˙9�:�Tr" <5�5���6(�'��xvM�w�
�����4�����h��_�Tp�"a�q�v ���[=ˋ]�b�y�q��b�&�׸�m��X(��W:�kbZ;�IT�k(�wl�PͻXo��'bH?�L���$��=���s�`�ݮ�Kx��{�^5�5��� ��d��?�w烡�"0u���W�	D�9�9# �*j+}��?�ih�rg��zx)ZlDeM����&�l�&t�'�)�O�{Mё��_C���Ӌ�s�F��g�Xt;��;��'��	jB���?��A]I9ՠ�{��żs�Z��=��>��7~�
���s����@�MĘV{V_�W���^Oj��/`H��� i���w& �R�%��:ң=�7�%	�O8�4�ֲ�YçD�=�	`�d�+�UR��v�S�����K�;z%���@���1�I��1K�A���[��
C��@���D�d��nO�����^��5�!�y�t[�T�@����laOQs~�!JBCм���K\���W������C�߯�a��݄*ڀ.̼�0� =�,V�)��E���$� YE���x$�L�"��
~�UT��:P�r�l��&��;	3�藈�G�_�{�/u`6G&����>���g�4�OeB�孠	o��K��,#Dz
R^^U^v����՜�|��I����U4j�u��x�p)�s{��v'���OY�.O[9O{��Rs�z^<��Ad�5_D��)��6ۙ����l<\���KS�/Ր�ݡ#Q8��H��F�H���N����]蜺@����`7)�mo�=m*;��sL}�`�d�d�Tp�rr��q��,bM�M�����bܡ��ֳ��_�ѡN�L����zX*���s�`xC}v;��%�R�[K��L�vl;j�\'V��H�t�����Ҭ��p}�_�ކ�Ms� �_YZ�9��]|��lYh����������*,c쁬�@|Z\�������֬CiΤU(�"�����L���owa�S��J��ڂIb݋���:��#��-��x�wg�ەw��֑�oՃ?�Ң��	͒!�jݲ?��d<�n�J�Xʕ_(҅�xm��>�и���J�z]`�~d[�eD�.���
P ��z2\�r b|��Q`o�����^àS_�������)�]'�\�Bq]J��&�m��1�#Z[)K�1��W�&��!�+���*��/X���8���5�� ���L��q�0�1/Dh6�!��O�kHf���p�uD+���=��eY�Ȑ	gؚ���y�m�iX�H�08W}��WI"*�<' 1{}��s�]f�Uň��qm��6����'O�2�_�<�W�vL45a��~��Ӧ>���o��M�����W"��AQej�k%B��S��@�T �N^�{����M���21�ͺ�)�Y�{P� A� �:|p�(N�3i!R�ڹ!]Npx�l s4}ޗ���)�I�dy�]�eL�\���ʖ�yaoD�b�kSB�,�'���I�Ab��v��������X�o�s�ꂶ��$�W�Њ$d�Z��M'�[J�� -,�O�i
��ı-l�r�>��값�<������]�f��r��MH���z(�����ݿ�U7�|#Ȅ����;ǙƻZ�4�lq]��c,�8�іhE0��{����X�|F�T�D����L�ވHE�w�w�p���t�n�q<�6BgT%�ݣ��(a��ٞ��곡u�]@��e��
H#I�v�
���A@��|�^.}ܪ'4�t��HrHs��L��,�2Dw��ć�.��������q0��=�3F��w>vρ5�ey���#ݹr �9�8�FA���+�f=ф���HU�K.��U\(LV��V:i��3�be1�O�:�Ž���2�Cz�����2®��n�i���l����[�ȣ�e�8�����]�Ub��i\L���l�zr�����ۼx���B>�U�Z�L��@Z�c���c!�b�`(��SUK�`5�6#�LX[pU��^������s���;n�@mg4�9��*|���ɥ6�`!����"��2c�G���u�}��Xu"#n*���Lc�qc4��+��n�܂󴢲(FT�;�1@U_y�mF9�ݩ�S袝��e�F�!����|U������' ���G��iv�6��#)��,�Խ����~!�����`�v�9je,;��pX�V���:x|�idX��iR���g~�*��5�Ee=&թ$_.��2���EY�0���[��JK�V�� j�g���_���"�4�|��RHԅH�~�t��f�*ұ�1d��9܉��uv����R�̔R`_~�� f���zϷ�4�NW���RP ��6�G�/"GXf��>	�2� Q���w�0���	�G@�+LNR	OcQ��Eo��{4 A)���uUEN:��+��,u�ma����鷤:���q뤐4�:!8g�:�⌒������~MIf�e�kS�u�$3�L�gO�ZD�φQ�E��>�Dx@��͆A#fk[	Ǥ��&��@�!� y�~���3G8���E�]c���>Ғ�ݜ����XQ	pH�(�dd�q�PZ������CF97C��|���l��y��xz���;�����D�nsi���a��PP��.������Q��~���f�M�b��G��@K'���w��@>w��^{�=9M���4������D9��W>���F��x-�� �Չ��`,C�D_�݂�x1�7�*�����0��D�K�#��P�ь�����΁f�uD�{�zg�-����F��;1B�c�),���Ն{M�$�S�t���V��}��(0��'H	���5����i;\�-��ڭc0�F���9�9�`����u���b�� .7�!�CA`�`c{�Q��R�@nќI��Z:���0��a��+��#��'c�g� ��	o�s�<�"k𻵪�)9�d+�������p��
��uj�>�iw�kQ��T�#�o�m�n
��#�c��a]㶉#~s��%�H����`x�k^/-T�=y������d:#:�����f�TK���id�F�2�Xv�w!��7���`e��O0��O�/�\���.�toq�eH�qB��BY��ŴJ}�x���Sʰ�v��\�އ��]�x���2Kc%�z����С��#)�G*����&^l Ő��C���:��=�QV	+��x
��BC3�C���⠱���n��pD������Is
���"��MN�[��c�	�!.Nߥ��,���sa��q��bhR� z.+�3^�{���<�܊3.�ܥ�~�Z���8��R�NHq��$ eg }�DX�@)��5�R�Z�P�dE�x�},C�8k}�3�:AT��>�kyv�p��p�(K�����������W�NQ�����q;��Y�BP ��Rx�*�B������7��p�h���H����F�?���t�dd���X9�����/���{ץ^~���;�B	�N�y�>��lV��Yf�iH��2���K�3_�o>0��1�A�a��bL�I'�Y�]9
�q|}k_���P�n��Ǘaƿ��r���?���lmj0�*�|�	F��8J#K�݅_TPz`2�S:�L���0A	12C�W�hRϷ�+O�U��1쉇Dr��}�E�mvc�rj��<����X�CxdG������Ǔ"�e�e.J�.���g��y�u�k=w,jI'�w��l�x��
f�˵0���S�*Z���"�8��i?����8��qw͟�cIÓ��L�B�c#�(�[�1�x�
���l�s�U�% �����c�y�0�?}&�s`KlYp���]���k�ܯ���kZǭ[z�*O���a5/]I��RN(Y�@d��SOΥ����G�aP�(Z�"ٸ�챶.׫�7�1�O[6��z�B��9���'�o-�M����7�>D\�?')ɀrp�孩��5���>,3#ϡ�t�i��6�T�Z��.�3i�*^(���� �Nt�wМ���G@��'�2u_>5@ �H�20��z�
<r_3�--Xk�sE�h"�V?�/�q����?��s;��}J�P��\���P�F� ֩̅)��Ruh����b�=�����b>�
�(�-�>���}��]��M�R��ݬn+f��3g�!����V��Nt�Nc�O~빱��K�z�¥S�0)��HD���t�S�T?5lJԥ=�U��?���ʴ�O��vZ�[c�����5�K}��9�ߊ$pD0p�6��>��[h]���XՇ���CJ�����Y~�)���(�l�`�e����v�=� p0n{��J`cfDЙ����9���lr��QH��¬ʸ~�l�9�^���s������ϓ/��@��闔�O���]������.0�Z2�q!����}�iW�����y��1�I.��Gt)v������i�F��ElF�
�}��~���3�E0Ƞ��d�q@?� �W���v�#�C%��b�K�ϲA�>uO�qnb�8�;�?��6S\\I����BV�u���WTvk��q�������j��QE}��E�kEkT{�*�M�'J��Ex�rfLߥ���x���Ϲak|8[Z ���7O2j���=�P�v���-ȣl(rZ1�z�6��+?�ğ�
�N7�B� ��a�2���R[X|��U�f�w���M���]+Y�~��xZ96�f[�y��_��<N�{7Z�c�lL�����L��Uk��7=�I��q�r)87+<�5P��YC|��}f<.#4m��eZPr���y��@ &Y�c'�_����0s�E���7�`���w�r=�w'���郘+�PlGo7r(�u�P�%;��c�����4�K��r��K��9^FLi� Z �
ko屛�cL81;����cv�&���隥���1�]8M7�gO 3�n�7o�iSȯ"�\p�KBHs0x]\6�a��4���,0~>����֣��e��ʇ5�@}��D�b�W��!�}