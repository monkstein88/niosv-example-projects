��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��0Ǟ���:�i�2����F��Cp�٧�%�VU��^�}���wWN#�|h2+2D7�ҸQ!��,;")E���A��j%�pI.y�Sn�ئ(]���Q�X�S&N��ߡ0������<�2��.�(`�b���ZTu���`�U'� �.�2=?�h��R���{p�mF[U��߰�ŔP��1t)�� �����+�@rB�ź,ʝ��%7��e��'��e�h�K&�NDِ��E��y]�%k��քچ���a�S�D&tǿ�j\��.�D�'eH[ͬ�i���i��&��TU �N���@�:v�Z4�{�D�B�G����������j^��=���~��bg���P��t�dn�����ښ���tj��Oicr�}H.M�Cu�X�:��0C��+ ��~��\f�")�+W�<��n�擵2�t�����5s��y�<fsW^�0|���{�yT~�c�R��R�H�o?���!w9��]1�Ƀ�]kv��E��V�����_~[��p�c��wj���#;���g	rc������4�CqT\H����肢����� �j�Ehc�D%�XH��'�:1��7�Lw�[H"1n
2�T����	�!,2S�5�SQfq�#Ȟ�(����( J���d��[�l��#��8���tsZؘ�r�V,Tv��Yb8��X��;ɪ����G�]6\t�ʹ������?V�F慑���u����h<�^N���� 1��������H%TN�C�ƅlN�y�=ʖ�[�~$���%Z^�p#�D�	o�L={,�͟��P���h ��G����&ɼk}0��ٶ@mƝ:�j�BBr2?KN�l��?�ǻ�9�E��F��X8���9tn.�!��V�D����Zx�:��	������F_��O��+�ijgr���ڍa�q�	l�/D�&.m���:�J�dCW
O����j]�%I����a�=�/
��@�N1ѡ[�ddˮ�����A#p.�$x TD�����t�WL0 ���*�F� "�1�ხNQ��[���D����@^��0$�x��LT�[G��W���	{|�GW�,d+�P��L⇵+́f�������6�������U�9*������Q~���\��tާ�lP\u^AVRb���:�� r9�]�?�x�J�꿎g<gr*�����	��p[���D/�5�D�;�b�}�KE�5��/�f!�eX+[��"�A1�4�6[A`��e%?�	,�'��d�`q�GE�F�%FA�׳�ր ,hȈ�!����%]|�L��1:hp�+(BJ���ө����]RG��! e�m���6�v���@	%�5�{����w�,�|�S���LuO�Ċ�6~H��K�C��*���dnW�͘刀�DL&���7 ��� ,�=v�c�̺u&1t�/�J��d�K���t9g�9�n�Z �!�/SA	��()�,�4����a�u�w{waJ�n�O���'�E�|�,zA]�$w%��y��:�RU��CK'������#`qX����`h�����N�ϭ]��p2y=�,O�Bܳ�A��Y���r��~GКw*���ɍ\��P�E�S������W+�-)\�8u[�!Ů�3�oES��Ὗ�<����Z����xr�0fp���R��@��q�0T����dPe��O�$b�}��/���;8;�~T�k$�M������3&�5>�,�G��� ;5b���e�p�ʆz�&ە��8��AO]���я��hT���4����O���?b$�F�9ml��[��|5>��>��o-��kK�ċ��#A��O4���;Ź������d,	�?���l-U6���yMT��bgt�B2ι����q�veUw+,��.���@1ktj�ez�q�����'Z`�j��=t}�e�-�������$;��(���+��=�z�Zx��G�A��E�بǮ�'{�h'��×¤�z�Q��_*�^���X��pS �7	$ڣ�|�>�jP9}x�!��2�=���Q"�Z�Q�E�8*�ݮ��.���c7n�Âme1d�&�;��ah�n��hb"����#pC�`F0������'t����@����X�_l��b��3�K�/F�������_h�Kw�c]s��{����He���JB,l�h/��`̲}��L���M��Nz���p5�ݐ��z	D��J��6+d�G!4�`@��dzg~�`�؍�DO,U.Sn�7$a/���N� �mŎ���/e���������B��JOD_��w�-2Oo)x��[/�pQ��v*���PI�B`�C�CG�8W�_)k�x�(��ʑC7sn�Ô�B��biu �%��^:s@6��H5��}�L�|J��+$�����4�Û�u`�Y� F�ݚ��kHڍd�ט���)���f- �O�o��-�'B&¿��^#��ڨ�I�uJ���'��(SR�'Q`x��79�ј	� �3�5u��UK���p��h��F�7���[d�[Â��c+ F8�t�l_�,�TZv�95�U��յy� ��8�H�������HU��`����] ���A�E�Ŋ�xmw�c�ӂv�&+���� ���$aR�A\}��14<+�'�c �o�H�q� x��7JX�8b��F�8�2�$u
���C�ױb���-|]6��R`�!M0Bb�=}ҩ���/�%��� ���v:�5&/����=�ve���nM1�(���wu��%{ÌЙ Yv�`� F��zV�>Zw���% %|�7���#'��Y����C�p�nQ����9�hZ@������U���|p���jK��[�ȘOE��n%r�X�È�Z
�6�������Ƒ?��$7���Q{l��R�l^��k�7����Q÷�%Z��Xo�m��F�"�L����6�������v�i�Y���,x����.(�QS��/��Ku�u�H��p�m��`c��W���B�!�}�j_V�zDX�C\|^�9w�/H��d���hrq��åp;������j*{Gt����ݾ ����n=���p�@�a���'�h��)*^�I��5�s�(5x� <�����	F��]d���m)Ml~j bQ��G���a�r�>��sq�p30i)��8���%}���4La��13�/���d�憏��ו�{��I���JH;�,򗍀��$�_���f�L�O��퇁3-��d��C�&.+uk�4HD��^�Hz�]�g��i��d��Q ��'�!�ϊWT�]�`T��ۦ����ז��� b�4�1Y��z��C�@�]��*Ĕm����W�j�Ƃ���z�S��c��wQ��h>�`���bp >�Q�U�&~��Z�F���}p�3��u��oc9����d� e��!�W�'���+cܿގuu��d���}p]&����<L��
I �Ι]V�@�"��Z.�%e�����HHtH\�wpo��f[dy�>���x9�h�,&gdj��`��Ⱥ���-C%��{a�O�Lպ2-쥀�}��ԣ��L�UR���z�;W��<B�#GQ�9��*=b�!7�7�l@�#����d���ҹ�,�OOء���?�ga���C~�#?;���]�c�@v�8��f�o�Zm6EOë�^�s%��+���Њ,���`�T'	�(^U�6�_!�#���]v�==J��HgmfaV��?�d�P'#�[+?v�񫂝t��^�9HNM
�V3��S�Z
�1͖=��$�'�NMܐ��-�Y�^CI�ji���1�R���7�ព�'e}�y6���km�"놑�Z5��X�Ti�0�ޓ��>R{`jŀ�P~�G��,�����E��ȿQ���Ϙ7�&����k��b�4�r4�	7J���&����_c"�+��������H��1�Iym�#������(���UrT-��5N-���3G4�T�ob��R�xX<�a�[�ZB1��~��H6�����MF�%R9G�O�ڶ�qU��ǆs^00&���:�A�CL��Q֣�p��L��Y]䓜�~�����=כ��V��*���L����������3�`_�	���ՀX2��eh���Ә�H�Y�//�4��2�b5�u�?]����mV��$tq������J71I�;u�M�OVd�M���Z��jA^U3W2���.��V�J��!y�]��2��ʾ$^܃�O�I�9��ρ�����>����}S�J-��s�0�u��G������1���8H�Tm5Է�=׃�o �����en�y�=�G�@f����dˉ�֨K�ϹE\� �cH(��M���= ]�����_���,U�w7dlbĲsF��)�9Bv�>Bz�4�&v��&I�-���a���| 	���(}4pVt���\�ufh�I��N��� Ɖ(_����tg�KxUt��<ʔ8���W!2�����W�*h'_Xo����uTכ�a�HpJ���y�Y��'���1���d���6������3%���adD�{Θ��@V��d9/ػ����I 
�)#\iW�/+�R�����}ξR�J���X���&T�����s��c�va��/��>tDl��v^:7~��R���K�&QS�>���������ҒGm{�4G�c����?���� ��B�!2U�n�������_��5jQ[�X�@�\� Wve��"<��t�˂��y%�$����7�"Q�HL���ݽ"&�e5X���Vd"��A~e�%bp�P�D��]O��~�6���B�8�t¿Wr5R��TVUX����t8\#�_�Q0�À>�=,�"J�{��:Ic��k1״��S�������z��%��Tn�8g����P��:Lw�f�s>_�c7�-��خeތC���g�	;A=d��-!(hp�uޑ�|e��v��N�l+j���J�CU�~
Z��BA��OUo�&��[�
��ިz��e�`�����QGPah*H��3G�Hr<DU�H�aX2��<��j��+CP�l�>e����j��~?�\���uȳC���Ӈ��<!W����{̀�R�z)LS{�PvZ��*��X��,����,��z�J�
�I��)��