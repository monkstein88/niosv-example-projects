��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2�}���i�|�>�C�I@K���,�>�����ȑI��)<P��,|w�4��5��Ij�$��	� daI�LWG��k����L��ɦ��6�K����өv��Ⳗ���	�3h���
'�ڑO4���0	�6Rw��fǃ�4�O)p�v�\+l�;�٣U����"�Zo�-p3�#�� ������S��H����f�9� apds-�]><z��]�H�������<�.?&8_}��f�Zo�� �ىx������=��Q��^c�v$�k�ڲ���q��(P�_@��;<�T�g ,����M�Iҳ,=��	�<�!�wD����L+Z�eB6��\EE�zC��BG�܄0n�~.c�V�:B9�+\Q���� �X��g�i�q�2���k��LPN�4�+�o��h<_`����I))ԱQA�[�+C8"'ɰ�~W�T�ˮ�f�g��Q8� ?K���4VHkBp3�ªg8���.I!kU|P��%����z�zu��}��r������e"�9M�`��ϴ�[d\1�>@�b����P���'k����؋̻�{�6}��փ\\��B�l�e�d��T©�;���}�k9����ދ�q�o�v�%kkB��n�:�X����D��g͖x�k)�Y�� GK�����{˸�a�M >��Vt�{�s.���S �Tѽ��1îV
�Ҏ�!��ɔh�����kȶO��`m�J��M���kH�w�x��U���x��D�_��*l-gl�?�F!��w8	�tm��8׊��g����!����gq��Ӹ.<2�kf&�%������F����$�Y�jqG"Zѐ;n���%����ߠR�x%�mJX�D4����S�1���KJ�zVH�|�DcH�{�KDb�&�m�VueZ��pS6MV���&��Py��p&�M�Xһ�g!��h� �ʶ�ן���:�����%#`aŞ�!�\����̩3�ގ���˷2T���鸰n��g+�9�S���\Ṋ��s��%*�%]CnW-x��d���B2�Z��V+$-�ŧc RU�f����qh��B:[���?^ꩦ�n	��=s?�?Þ90���I<�g���)�I�g�����I����8cS�W���V�]QYΏ�Il;�����x�L`܁���I7"5�$���k��b��I�/�ŀ���@E� 潷�q�^2���� �ǟ��6%��H1&v�d�y�L"�|°I��*G���
_�_�DG��JC..z@���&�(�v�`U>fn�)��JBDn%�����q�m��ċ�Z)v�.��
{�[��+t�[[�/s�lT�u�^�T8�-���g9�����8�#x�"?eZ��
��ʴ�1�2�,��O�h3�I�4I��ՠ"_f;ڒ8G,�B0g�,AH˜�_|�!���7�6��W��෸��{C�d .E��)WM�u���3a�+3J�3N�)2%)���m:�
���=�%��̯vʩl%�~3�ަ5w|�� �h%��Lo��A̭]+�X2���$\�e?�)Q�iuݛg-lyaHKJ0�w�b@i2�Q��� ���cֳi�2�0՜xG���,�ƪ����q�(
��ԍ�rYH$>=t�:�5��>�i��I��z�D��S��p]&B�YN-da����k���Mh�@CdJ�mJ9؀0O�-c� 吝
T撌@ZWҵh�&���J��� :���@��MFh��G���DqQE�:�%�Yk��Ƀ*��P�����"�w"phI�޵�2|<]N��Z;3��tz�E9�i�<��\���� ���B�B��\��I��Ś�����X�\}t��gd<�>F�GR�di�N�m�Ư�ud�{\8�w���� ���ߢR��� Z�R̕q���3���M���e�����������s��5�4|o�c�N�#Vq�f�}S��Q�eg�k`���o6�)!���~&������Rny4��>MMq���0����O�Y8w?�� ��Z�i�@F}��ݬ�Kꂣf��9�n�},S?)���lP�w2q3��?��\e���-�����*�|�f��ġg���A�dqa��:� ��d��������~��(��	Q�7?Z-�5�J���o��~��eP��+�7��M��iEEO �����Q����$����ԝ�4v�笢уѥ��R�����_ �h]�5���V��Ʈ%���X�H��^>0.T����s���<��A�Q�80�=a��`p"#Ss0E�=��>����|s��G��p�ݕ���x��n�Q���[V`�0��_;�p�0#��1��0-�O3�Wl��l���k����� c$q/�<X����2}v�w���{2���o����1�yg$a$S6}�yQT�X���68�r�c�X��B�����xNDk�t{��U]� ��`=���-ޮ &`4�{�R�j�Tm2��I ���L�=���)����a��b��d&�����I�ig���h`sw��@/���H��(����,�G,lUV��(�cj���ոƕ�ԯ��u���x߮[���L`�wx��"� _��4>���U��"��u
��q��]��ª̦�|��7?S�g��0��G^���w�'-�x��[��cw�O��0���D�l�������t>+���ԯ��v�T�=MD�ES���2|�3=i��պ$���8b��/9?%�e26��xr��5�"R	Hd��/2&e���"5ڬx�R5^�� R�i�Q ���b^I2�����-�cU�j��+��{��e�� �M�&�ɍ&g�{�������ֿ��M$�y��ʑP"'�a���r��5���(��MG�>���h\ !�H�5xJY���k1|��'z���V�k��$Q.^ܰ�DF2�7��nW�'���ʪS8 ,Q�
t�P�Y,���7��ܡ��h����yE�6���5��e�0.��~�pH��4���V����#*��	D5�T����\[����hW��_��q�W�d������P ��y,c��
~(M��VE�/bʋ�J^�O�tB9O��Sd�����3
�u����:��&y4a6ks_f}4PeΑs��(��
�J�޺�:��,}L�7K�.�j���g_%�8����r�������Eq�+�ކ�` ����D}5�������tf�	���}�]�O�$�L�*�1-vg� �nW�e��{������<���7ޖ�1��X��H��p�oj�)X f��r��CUƎ���Ο�%~�*�(�iDa����(�a���\��/�b�vЛ�ǥUgW%)��t�Xjܗ�ײ ���s����r���K'lw�� :�&Z�����2�)ǋڀK�R��o!�h��b�
0�r}S��*Si�>�{yޣ.����3�o{̥Ł�Otp�J9O_�J.$�ILu�mH���
l��NZ#J�{/�(Q&�F��v��*3~Xw.z46�3��x�^����Z��e�4k����د@�K���F4��ɍ�5f�e6��,@/H���L�ƫ�b��]���9���vQDB}$o����n$4��dn�q(���������Y���{X�r֒�>�N&��d�r���x?�=:���P��O����%�Q��E�в@^��4���Ñ��ߏ�Օ�uf��4�s�@PE���A���mm�s�W�K��<5l�ӜO���b���)�8�����}�T�֑��9�Б8�q�Ie0�G�h�L�í��'��2�uy��u4�wS�·�"'�N���jB,VγYĈ:�·� ��pO�C+d`[�
��Fc�(\�w�W��+M��j߉7���$���}�K�}"茄\�*��@TjBa��pF
�tD��0qƨ��:���[N��}fĤ��$��|������v�-�|
+���O��0|��s<4'?4�)-2���̈́ۀ0,�o(돽t��%Co�^�xwz�~�:)������jP�ʱ[Y6ЀC+Y��>�ƶI�r*��9�c�˩��|`$#�>�z�b�E^k�����st3+EyO�nys�aj���,n�ŷ�t]bRr^���b5	1bnW6j&��y�CQ�"��j^X���7�{T ��n��O���q488����md�#���,�C=���p��8�ah8R�0 Hјq`Ms���k?����:7$t��gh>�� ���>�^����Յ�H/�#N4�X��
 )��G��f��Dv�u��� w��6�x^x�p�4��n���M�_�)��(��a;�e>Fs�?�h��w���=~<��Vٲ c)�L���p�uK�7�7��p�VZ|=�Մ?fW��P{��g��y��9����D�o�Cj���(�R"[_�Y�${�^������Q���6�Аs|�^��w�;�-;7�u���|qVR���wo��:����4��P�%��6Q�9��H@S	@���ż�l/�w�t��.���Hw������{��Ĳ� @�>Q���k�{�vf�$��2D����;T�k*��wuH_8'x��m?��G�YLM���2��<���F�M]����a��v�����-7�kW�.ĵ8׸w��a�����	?U�5�O5?�o�ä�ߡ�R��S�G���'���el,U�)T׍�`��t�R,XI)J��tnx1�i��-&Y�[����06|%�%+s������U��5w�˔7[���Ԉ�b�'x���;])������*�@�W��/Y����Dg^S�����Mx�ɃF��Y�=��H�`�����`|r���;g���U��T"�0.���2IF_��C�����A��4^�9�d�O��3D���q��^�B���.���E�3��Kh�bLz��X��kBdfb���?K߮k"�/�0����x��
(땮5_����r��\s��s�ޱR�$�o�� �W���J��a})k���W���
z˾�_n��W�x�/TR�op_�� ���*����t4Y@��U!��^,�:]
G�<�m45F�J�`���Zx_!�3y��t�62B�܏�a� y���@���fD.�G��q����A ����C 8�"��}�-��ZJck�a����e�9p�gsӡ^a}뚠8U@��7�}�6��_�! �o!����e��ٿ$A�
Mb��J;��N�X쀭�S
��Un� ���Fx��Wm	��s�Z�.WJ\QE��,�k��픳&��O�p�p�
�t���*�{���T�� E��ٖǣ��3`�ϺN��慒h��mP� \���ߵ�n6Fd���z����$A��P6kơ�7P\Ƈgn��t���*��fh)��&v�ǥm�,��pB<-�C�	 YeJ3���o3T�@��F*�����F�q��-�cCmYP�=9:CW)�?In�����hH�y\��6�]�\�����;%L��m��݀��k�1C<��G�f	��~M�/&O�#�� �Z�k�M�[�^M���pp��p�8`�AJ���:�/���Xuqͳ8�r��S��|������ >2T��o�9|����y�
��W���vbp�ޫ��%�"�Kt#Q�
z}1�pZ"6��	d���:���O'��kț�,	���_�5ԙ�sH���L7�(Es��xrʛ������e����)F���d�r�g[3��G�P�� �raL�t��o���v��i*�@�Ę�x��t6c�� x�Ӵ腄RZ.m'�/�@���2|l!��񎺅M̙7�yB_&��G}R=��g�D���T�1Q�xN��W�U��d3�vZU�Vߞ����9���z��\�|<��(dև�� �pZ[�D�Vodj��<�%1a]��ݒI�s!������_����X�>DA�YjV�uL��-oq��X`�oM�MN�~r"�+S�ז6pBՏ�mu�6��IQک��>�@�{X��b��2	��W{���d���R��ڮ
u���	�N颂(8OÃ"�S���R�p]�8�V�Yo%,����I��mE���\��_�g8M=�IR·|E��Ԗ�H��Z���OP�:�'!� ̲�1���(�+E��π�3�%iB�f?��>��b
 ܶ!�$w����"	��Ӡ��P�$q�1��@�u�;~�/��U����^�3�vS��L��. 6D�Җ�rg�h�o(p�m��(��}���E}E����u5��6�a��V�6�i6bH<�ū%S~�|n�_��\T嗤�'���wRs1@ p%:E��y�{�y�Ҫ��!�X4d���D��J�Om�ZڒX�tZFL�{)�fѽ��j�s[k����b���Mǚ"����ݏ��:�w�ć�����sx\��>}G����W��/e�z
V�� ��ʣlB��O�;�HA1�kG�ˌ��H���U)J�፟B����l����\����jk�p)Rh

�]�U�_�Ju���������+��~;��O�C�w��}�CY�|C*�M�+jx8I!�(���(r�[�,�!Dt%i1֐Ad��<����q����('�@�w�Kx�[<����`MC)���	
��	ю��Ʌ��X��(�)������sW$z����^��3��QA�p�5f�-p��"�R���e;檂��0�9�\ґ�cbq�>D�<.�K�����m6k37�G���N����[-[� Vt?�y�����W�b"���H��a_�l&@[�`êz�^/�?g��T�%��uB��y�\(�.��}�1�`�[�J�aG�^b>q@
uʤe^,���̂��4�H���rK�$�Ż�#��$a��/3H��VC��Ǆ6��W�VY���a}U��h>BZjq�$�V�������3����\�tN����xǶ3��A4r��âJ\���LG߇�Y�}�^��j�����>�g�3G�q��ݓ?3�E��m��2Pf�D�j�U�U(Mq^Y�h���<[�3#\r3G/g֎+�����"Y�`�2�)9�H����+�����ߕH�@�����9��N\�wUG݊l��u�!N��`�Z���� |�U���\�#��W[X��!\pm�py��=r���8X�����Џ$���F����YU��7K���JzҔ�у�~E\AU�N*S>�ޜ�}.���o> ˒��V~]�E��5�a�\$t�r��loT?�Yzˁ�_n��/U�g� ����U:3V�7��rX/e{C���Dsܺ]pMpم��bͭp셜���I�
�Wޖ� �v�)�Rk�12T�m�˕�z�t�n���"�?ݑ���;��I�`����i�n��O}����Sӌ��)�P��� ��م�|c��Bf��w�#r�RL���%[��*?ֿ�2���&�+���8�����4�dWO��ʄ�S�E�^|B� �D�>�A�^r*��! �V�y䘤��TL����\N��9�K��
Ɖ�G�k����f�-��dE,��{��t�'�D��1�ٯ.%�B�W�ϑs�+x��?{��pv�#�u�~��
cD���Ђ*���2��w��U�w��-8�:����Z�Տ�ɺӵF�q}"�wM�a��l�c�4��]�o�p?�$;�τ���B����X9T�S����:���G��d�WyR{sx@]Qe	�!��g �p���j�O�h�4P�<����R�����Fy7¤+���s�:�m�nfn���S����B����F%W����v4E�]-�_ ^tn������4qA3�qU��5g�h�{�����k/��^GT�`�a^��+=9�Z;�;���.2;����f���J:���/f6OT�ٝ;�2hrVbb)cH�ac;xW�&d�0`Y:��?l>�.�
��@���p4�:��Y"���S��A4u�w+-63p��/��'��1`�=�xj_���T7!q%�0��lJiԙk�7�_�$Z����E��X�̀�!���%�B��9��K�D�S��K�r����74(^6?��q�Y�	��`�e+�;$�=�	����:J�+���=&{�[��S��J��ʷ�ݕ��I�D�Q���M�f�����J?�f3��uM�r�L��������sn���k�"�D]Ѭ%���/�`ziǗb���n>߳­
َ��٘6IB⳼�k	�'Nΐ��c�4S\<�\D`��T�F���W֥���+�#�1�i4K���ì��&�rvbcvM&���J�W���f~��z��ԮO��n��FU�����E�׍B��-�Y�+�r~���#㥖r�5E�C�T���c��V[���b*��!z(~U֏��l5M��j|�_E�Aқ�0��(7n�=���4�*=�W�=@��7�c�l�����= ꪍ%�ㅬ�T�
` [����X�Q2��K[@��`j@�A�t0�K%�}_<
����m%���ԁ�&��Iv�x��B�K󮾤� ��h���%tx���n柦����(�g�zH�?T�E�	UM<o:0��63�$�)oȮ�0�b�Β���/v��;2���VX/�ʐ�gGq$�\7���sl��yWJ�B(��S_��d�K�.�T�}�ɭ�ʉ򙥙���P��s�����>e�w�����Q@���z�'��S��Έm�"�&�.�|� �2?d�$ɑ�	FԖ��p���0��9�5�)����w�M����v���0�q���Z²��O��8�M�
���*y{hP�f�>�*s]
�C��-�B�ص�&��/�1�8�>���+�E�t.�K�Tu���(R�eF`�NH��1/��r�e���t��σ�� A��΀�BO4�=��-�*sD�胭/\C���[b�OEx���d3ɂ%�;�<g㨋�+�s�e@q�߷�i���f�w5�UH+#��h�=ZB��H}��o����+�'��b����tQźHO1!���[Y^�f�X�+���D�T$�?Υ����ym�]���5G<���Ub�2�h����ⱀ`r��V.NbK�?5��a?@��$�e�������?@+ �v�L��i�Dh��(,��Y.e��7��%9`����3�SLv"݋*��G�C�K��j�$C�%Y���4x�勸�P<�~\ܐ�SxyP�E��I�ƥ���p��w9��U/H�Y�h�#:t*�{i$Π=���֕�������TI��UnO>  ��~�� s�%������۱�t���I��;��u�f"2.��_���>`|�Ͽ�~�S�/e��l�3愝#lH����l�>- @Xec�j���c}�+G�RY��8_����k`I����\z_�JW�]b��9@��;���X��t�+1�����.Ԡ�=i�V�s�n	��LO��~�M�JX�7��s��W�U-������|�4!��={��HK�"�k)�F8j?�<Ao3* �-w����iN��(tlH��jR:27� 8ɫWl�EX�[i�� ��~�Rp�-�qɁ�ʄ� ڌ�����/y1���]ћ�ۭ+��ٞ�r�P�`��q� ���d~�T��MZ��It�z�Yg�8U/0�~l��]1q�Sی�+/�$;���F�@Y%�Wk<��ZȰ޾��N/,�+��da��	��Ò��۴9��L�1Xy%-ӄn��We�U����`~I�;��Y�\�i�j'U��)_�!r�iב��J��Te4����Wu��ّ�*ۻ^4A��рt~ܺ�SÚ�Ӕ���TI1�r�E�?���_�P=c�e\�;/\�s�%h�2}$���%$ҷ�v����$4�94/�>^�3<G׏�+�~t�c{��/tc����c�B㷇�.r̶��orkN�5I*��e�Ӭ�V�/�ƵK�^JH���K�1"�{r�&��Ă	2.Q�E�,�B�p�_�?�һ�&06�y��<�s�˂A����v@����2��Ce��#''G9u<s��j]�|Y��o�l��-�M�Ne�-���e�3�|� ;蛂�ߋ�Q�:��>��R{Ԩ�����Z#�<w��ㄮ�2$�c���G~|%@qcCkK�7��`
|nJ��/��OO�LҔ.�Ó.!}�����'2k��1��WK�چױf��b@Y!���3�w:�e����wn��ֱ{F8�`�|?��Yך���	��批��ic}B<A�s}�0�8����Mw�N�)�*7|��J����\Z@�K�P�)?�"�M����鲐���-i�[@��VL6n-U�eZ�'3$ �!��&�=�7�=?�+"_�d����e��>nQA����8�ܟ~/y�3�2;J���eW�'�_I͸���X /�k��ˇ�c��}�����$���׬��0���D��#��\�&Gҟ0p2ǅ��&K�s��rTw��=ġ�Ո
��F�0�P���f�J�~i�Au��dR,��4�d��/��b4x��<�A�����M0"�Pi�}hm���j�`fv �Q�J�⺿��r�ZH�0e�����TLې�U?����U�a�4~u���� �j�uYԐ/h�c�B�=���mSҗV�K^�
�aʱ���$�2H�J���-�jOr܆��m6�V�+C�d1��A��a��D�F�����-�d����5]�O�"���0���b�Mgx�k˾Ҽ����<"��W����!���3]+V�A�u#����1�?�;*h�#q��"\G k˷�i�}е�VE�.l+~�{�ܙ.�#|7��=�ȯ��6��>Ȧc��C8��Ėm�e�i�w*d���?����a"��ǌj�đGZT�v��v(J�Ԩ��	�z>�ZM���/nk���������򖔬�ʝ�������g��J7y:�q��d����1�BI-PE�{ǌ*��#��ܵ��{�L�i�m�:@$+�I��Ks�WGn��*��t#�J��U ���Ra�:�k"��A���lX�Di�QhO=��LðZ�J�*�3��Ȅ=z�x�׎��h�C�*ZX�g�+�����!�X$眎k�F�B=~r7=�D���pFI��I����0���H��/1��4zit<u�sx��ͣ�V-��,�u�u�>y�%`�2�<s�=��0y����ރ��Gѥf���4�O���/����%С	С��	z��ß�ƚ�[�Ζ�^�C�N�nƔ�C	m���Fˢ��NBA��1���c�8�M��7�x���]�:Y�=+�9?��͑�3���)�B��t^�`����$��}���߹��2���A�7Dl�����h���s�nV���L�[$�v ��*������nx��AR\��Yz��q�cg����]����t�SԳA�R��-3�HR�g�MS��љVs� ��� ��6:c.k�/�4'��V���~����u�$�A_�6Q5 �&���J��3�ݑ�Z���Ǉ��F�����d�D����v�X������v�W��r{��P�k?��W���j�NrR�- �w�C��K����~�Dס��p��������䐕Ƨ[BG��g��'��kco<G+r��h����W�Uq�r���*ڍK2�����厍0�����UT-�Ih��։,���
�7�|��B/�s$o��o�>M�?o�����F�"���llb��n��:m�' ��O��1u�	�w ���@�K�F�t��{���-d�xՈ��j8���Wc��Rmw9Ֆ6���Ү�i�Ys�׽V�����\���B��l�D�\�cÐ�eNígM�/W�n9㝠ҙıWm��a��@!�w!(���ka�䫩�b�`�>]X~�U�ڠh�(fP"�5�g�r�,b�m�]ʹ�aֵt�`|�2z1qST�͍.�\z]Z����h�u���G��8ݙ�vH������\l:�cs��D�e��qn���P�< ���6>��m��'���%fT�6�"ea������S-��3�����8�=��LV�~�͡7��0�P'<,��ʑw��G�ڊþ�A����Bع�C��OM�a0�r'�JH�v�5�I�} ��S��j}g�d^��b�ə����k �1�l3���E���cz�4��>�\�
�dܨڢ�4�?���=̷�6��<ǒ��x��K�?[�m�,dP�U� ��&dW���?pXP�)I�vО��� X�x�G���ȶ�!�,�A��	n���"��U�y"'��0H�͙��l_���A�,w�4�Ȳ�&N���m�|��s��fB�4��cD��3N�^��"�ٕ�)��L/p�sm'�������%��V��R.�3k�?,m��g���:�Wźɐ�vc��m@0�3�G�\�f�p�Z^A� vV�[��A�2R�쟳揽�W����g2-]*Đ��!s��H7�3>E��s�!�V� I��#��D�D\��g����?���� ��"��r�ϰ^��H�2�8A{"������0<";<&#!��"��F�*��]f�&Y{:����IN ��^pi��q�k],@:��hS���f7;�'�9������MD��D���������Ys�7x���Z�o��|B[I������j�?�,��:�ݜ7�{�����Ь����Nb/B���Tșh��V���-q��b�5gN�q�jfi®����W^�y���Ԩy��δ�]54T�y���3]"p�O��0f���Yu�r��>���.��G��)QI�����A�W���Xl*�~�M���Ԛ���U��*�
�'��$RfM{�&O@��Ud���<�ֵ���>ҩ`��YS��M�s/w-���B���e%8�쟙������b��R��{��	uk���(�ۍ���<?94�	X1�Ϝ�����a;_앀���1/���>��y>W���Y�w�]�:��=(�s����SA�c���$k��ň��wERէ�-BId�P�2d5� ��37բ]R~Դ�[L�q��A�1PH�-�֫���,�72`���AxG���}�b�m�a����hL����ج:O�7�	5�q�Ƨt��y��E�����QY����X�	������ �>oGB�F��	m��y������X���;�,�Ԟ՛0R ���>7�n����A���rP�� 2���pZ��3[�w�W]��Tkr��@(�����bb:X#V8���<�Q��Y!��.�u��<��M�n�i6,¸�l��ˮh��f�@�4�@@C��rg�)DM�Y�{ۦ}�Kz	�C 
V�>��É��q-
�S>��$�N��� �i��?�yT�x��_�"瞁�d�4)�Ȭ�I�׿xe�|�e�-�D��I_<�8,��X���"jA:��v��u��N���,<-^�\�T^�_�}`�5�=iQoK�^Č \���CR\J����Y_gkk�a��0U K%"�i��c��31F4*���!� ��r����sΩM�‭V&-�0��=��/W�;`��T�`|�E��u���SǶr�@8�צlW��QUcO��P��L��p ��5�ȹ�H�J
��B$4��V;M��ϕV�s�jd}��x�.�oC`�5	:FG���rFM9 �9B�Z"�ÜA��h�ԯha1۟v��$��y�?���|AC�3"�^�G�`��?�yg<Ԓ�����n~�y(��>�b���Ep�l�a���3DʿE.���&�Q��f4��L��es�Zl�-�步���a��ԍ�
J�=�wGH0`}��.e�Q�>A���T��7=k 먷�^wcv�8nZ�7:�'���LJ���gݜ�r�zw|S�9~ۛۇ��d�В�F6ʟ
��R)�ox"����A�N�$�s'�7���n	�-as��E�I���p�V���Uh��Y�F��t�C� ���C� ~|�siP٢��'��;��G��er���$z`j�hJ�������n�Y��z�:'����v��u-](o��V��0(���}�o��1a�А~�ۗԇ%@�J�4%̀8K�����c��M;�d[jc.��U�ttwx��xQ7��c7)�^y�'�#��e��R��K� ���y���-�2�e(�y8h�(L'X��� q�����g8���?�t!f=^F՝R#u|%��� �qz�A��ٻ��U�k�Q�߉74i��; ?)�8��3�iY���6�����]����du�D��1���שL5�]@�vD����Z������dQo+�x�&T�v��~ͧ����\�8>eu��]�i^��������+tOdƹR�]$ʠ(]Îh��CV��R�0������=F	D�絗@I�"~��œ9Vsվ|f�eU�h���\56�d�C%�_@�I�<��dn��!k�؛Y���f�"��Y�~��<y:ݗn!���UY���<��1h�D�52<^+﫞d��q���������|�׽�����p�F�E�|�8fՙl����?mw=��e��ȿ��F����5& �9���ax�K�F����K}�̊C�܋d�|a�a�L���v��_S��]�{Vo p+�T�w� {E_:;y�"�"�;�S�0�I�2��|%VxU]jI���j�(���2�ձ��)����W̠�Sq�j�9"b��0�ĸm�k�p��G�>[�'Cw�߀t%�z�k�@��,�+�2s$�	�r�ZF[l��=�N���F`^)��_��D�0[c� gG5��z�9��B�W�1`a/�2^6�|��dR�U ��c��~~�F[�Ԡ��ħ�6؈�bdK3M,~̢n�VʞO�v@S�b��Ci�6��W��x�' �$$>�p�f���5�K�(��)�7,�	=��5�b:o��B�P�]�dn�0��{��x�xS�4;Z�a���-���Y��~8����7h�� �����*w�ߋ�E��c%d/�jS���%^_R�K3����(0}�*1,	,��� f�������ǝA���_����1�l�D4��x�� ^Xu� �ˏh�l�1��q$ �������=S�颂?#�D�+X�]7Z�)T"&�"7�եE`F��8`R��^֐uU�$H��B�J��3���D^L��Ki�Ϝ��y<P�jY�q3��i��5>��d�C��_�%fx7����Ŝ�֠��������%ީo9xx���?�O9.S(�~S�҅�	��7�ڕ���i�g���W#iJ1�y=��U�gd����*m�es�����O:�1���-}ޫgk�r�^�J����C��
H����v���"���4�US^9��γ�	K���|gۘ3��E����<�.�YCMs�+� ���q%r��$�0�1c�oa$9k{}����q\W���D|�S���N����N�a��!��c������:{r��A%<U,�>�rv���NEtjO�˫-O�����7d�"����G�R�2����a8����x�����'�e���]m�y�Kbq�����j�~��x�*S��>�6����`����1�=�WR>�0r/�- r�������,K�1�7�ބ���ݏ�j���Y%Q��D�<���?�����|������*5�����`B��ݘ�H�hm͠�f���x���d��=�O5�G����"��J� ���'w�zT�cYug��͐��;"0t32�z��B'��i���˰��[�Bl{z���B�h�'C¼��e02c�5� ��jl��*(��j�m�
��<io��)�(�cn��-�%�.��S-��	�nv L��������\��g/M�d�rt��2�IL�Y$�l� s�M���h:D�M87�՘#i4��GlO��	*�.�,wNBq�)�;/ԃB~`���˪2��R�����[O۸�U�~�mr�n�����`�O�;ꭐb��E�+��6r���N)$w�u���^����ǍQ9����d>`��3 s�ڶT�pkcc�h�� j��	�r+�R���é���q����9���o$r�8���5�[��<��ge�/���1�O����-ʴ`@�2:��IB�Ei���]�ޕF�_W\��3r�T�i�ܓy�	 �G<��g��
_i�ڷc|Ȕs4#���ߍϪ_=�&�Hu߲{�:�D�ˀ=��CO����֓y�R>�������XJ���Y"4i�ɡ�p�6��ēt���0t�j��:�Pϴz�_�h����Ũf���9'�kg�� ����-.�F����j�������R���AlKԳ���x�|��T��/;�����6��f���7�|��%V'	�ŕ}����=��[�O͜�^/�z59Rn~��qҭ�N�gx[�LiWZ�^%�L����d_}���}uN�?]�ʁ����h��2}�=�g�KW��BL���l��0+��q=+�d
i��ʸ�1m5;�DS�m���b6���nZp	ܭ�Co%�j#;��Z]�|)�}1�d!��,�x�I���(=>HZ"�7ՓZ;%�����]�(Xi����}�;M�{6I��9��ϥX|l�bq��=i��@)<G9��ܵ��Ēz�k'�$܌*��/qX�= ,���B��G"��k��m��<p��Hzu�V�&�<|`M������Mc'�Px\Ԭ���j��}f*���٩z�[B 8�y��_�4��z��U�H�x� !���m��+qL��\�І�@q�T�e�7r��u�"
`��z�z�:Am��Wɞ�n,�,���=	>�X�?�o�׬(5�WS�y�&dߧo�!��p���B��>�����D�^�Ao��u��Pg��JV&(�	NCp�hܪ��;e�-�y�ވn�v�k�Ǌ�[�9O �D��e\��q��N����|���at�����3l�G�ELh�$�� ٟ��H�~�	ܑe�����=�<�� �Z��w�1�Q������>u!Z�*bF�Kn�j����Ȅ���Xg'��t�a>]~e�QʪnWr�7���$뾇k�N�!�����z����n8ɔ��3|Ul���)���i�˴��
���s���K����]�+z�B�9�+�FZ+)H{��gf�Ծ���0����0�;ϓb�6S�
}�v'|�P��$ԪW@��k���bj��4�c�4�U7�6�KNH�m�Mr�!�0�D(�	�p��ҙ_Y8�o�KU�%��{�(ǡ���[�3R w�r���+�#�Ŵk<���]�H�L��k�k�Xl�6�|��V��,9�]G�}���D&q��� p��˯h-�>G�F�&,P>����U��=c}��va���#�	u�O����PQ�B��I<4� �#:�{�f�(�9�[OP�C'T۫}����J>�/��ag���ɤN5zu�N2ԥ�	n�;4$e[M,t�a�Cq<�?�B ��7B�$k���m�	�^(�A�]{�1�;M��Π�ʹ����wgG#<��zN�:�)^�2�h�x�:�7~m�y��]�of���Iߟ"�s�䋳�W��ax�9�B;Xy���6��$�)�V	����R�C�T@}N�p������z���ޟ� ���&ѿ<�����x���|`�{�ǘ�V�N��z���Y&�{�:�,�c��/�[;�qR��ֳ�[
�B)�����<�!��󏩮i�ʼ|)c۷��8nB�	�eXI��I�'L�,at�2}�^��8�l�&7R`PB��Yw_��@aVє�����=�����B�QxL@	0��!��C��<]�����U�R$]]�cqh����C_̴�_�}� 0b�������c�U1���v��سf���טy��Ed+o���.�y�3����J,�;[4�$���.f�q_>a��&=�e�l/�/�8��f
Ue	2����S��]vʺ�=�~��I�c}'%HQ��
~�b_��������*���K\��K�ۈ�E�d$n���'G_�6'm���w�W�kK����m:���d�zQ)<SΒh���;����10��Gt�o�㦝dJ�j�̓(��C�`3A��e����ޖF���ID�|w��:��q�\�k 暄G�y{��a|�W���h�Ԥp��4�B~v���tڍ#[��|"��-��l�c���(Rؘ]$T�Eb�|�����ۂ'	Ⱦ��!��@G��u��"=��D�e�wv8�/��t>�y[��z3������A�D��@�D2y�t�����~�Pea�Kր1�x�A؝���L̡x��v;:G�C�J�*ف�Z?S%�ֿ,�	�aU��k�S�cD{M����=E���6�x_׃�ތ��AI�+*"G���6
ߌ�>�֭པ������`%!��Ă�8�$��.��&��	��õ�{O�H>1ce3�o+�a���s<���ӧ��"Ŷ��������.��]<��y��46�r�0Si�.A��$��r�|\j�i"�3 x�ؓ��Q�A�^,�#�8c�	wY���y�I�bc�?_޺vw�!��&��U�����m?q�����F	hn#�g'��w��9�8u���G Q�A�!���0� �/�X�4lj@�Ƈ��� �چ.h��X�u\-c��
Y�<��}#tAW��B���2�������]�P$�V
���T���yQ��彀xkW@�@�Gp��L���?�J����S�E�����ƎR+�.'�:0���^��ݱ4 +J�N|�=��,���Bׅ�M��*)�t�٢�9��A���Haf1A㌬-�[�A~�j�:�>7]̏@2�U���Ft!�K�?`t�i﷾Ϛ4R��n�S�i�~-M���5~΍�n/�wvV��g���tիI����狃I֔3�g#e�3��R-���g�l��;����'���nY�{��079�����1`1�ωܘ�&����ީ'��=��č�/�L{����͑t|����DRu�3<�~ձ1B^ع����3̨R�[E��N\s�Gl�d�Nߡk��������83[�8YkoV~���(Q�0��wO$�uР�a���$�5E�5��N]n�Ux��MO�G:��r*���L ��1�t��}�ъA���B�Q�ʪ� Y�$�Cw|-N+�ׇR�g�Ѧ=1"��-��8� Aq;�騭�FzE5��@r��܍��=�=�/�B0���3�ôR1f&�-��ۛ#��Nhzʘ��p3(���7k��k��źϕ�{�R�YyY��]ܳ�c[.�ݞ��N��tZ�n晻�G��*~�2�?{lģ���w��'���UvN�� ���