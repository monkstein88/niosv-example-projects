��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��0Ǟ���:�i�2����F��Cp�٧�%�VU��^�}���wWN#�|h2+2D7�ҸQ!��,����ץ��k[��?B�����p��O���m��(�t���}�����P�<T���(�TԊvrx��H��$��}���:G�`����U�{��y���xn�c7;s��,������qڼ��M�����o�2��	_?8�\����zߺ�֤�={G�	�.0++x|��;���!b���$�ee���b>����۵M��9��<9����ʗR�կ)QT��Z�F�Nt�y�ފ�D�6J	�{����,��C�(\;�i��d��|�R�-��<9�0w;�#�v��	ά�7��Of���I\єJ��7���i��`���o��ܚ�K*��6L���+Q����;N����a���{�I��"�W���%��r�C1~����Ȭ:b ݏ����܅:M�0�F��"C��U��k}6��[ࢗ�\]��Z|��$�8�;�W�r���+f�%�/b�4R��:c�A�:S�����T(�@$��e��g�����;�D<���mٮm�{ f
��η
��G*�a�;��S��,a�;��Ȁ"�A��"bD�3o:��W�H��˹�T�欆yd��bP�����w��8wv�q�»MJ¨N
�O�&\����Aն�
vC��|��N
S�MN h���wz���ԧ��Ψ�-�[H��y�tF��!��glK8N�`��j��y�C��}�P����f�9V��DO���?#s������ƀo��R�7o����+�-p	�B�Eoq��۾k�6O�cv����\���>��h���6i���:sԦh0�]d{��]GБƷ�98Q�~��1Ni��79-s�C�4bm�<���^ii7=����x̓Eb�3�a.���������!Q��{�x!H����,\YUW�qmsE�ZĘ�@��_Ö��뀋f�Ddbn�͎���N�������k	���Oh�Q�������:	*B�L�"(�Y@y~�1�v'Ţ(ݶfޅR��x���r_�+x�:�T�O{N������2�-���nF~�$Z��d��7Cy�K��g�eU�4m��S�����z;��}��Y1]���LB��|�}|��v�M�>�X�$!)�z�or9��N�i�n]R��6�vJ����t�\4z	����?M��'jc�p7�S8��\�ĵ��+�'���ktQ&��U<�;��<+���Qc�~�����$Ļ��Ql��\�_�Y���K~�a��(1%f]ةdJ���Ss��`�>i��#�C��k��ӹ��k��y?�׾~�%���S��,ׄ$�w$k�h]����֋{~�W�~�y}�CJ��xq���pA��/<�ύYZq1�d=)h�A˵���oP.���ƾ�V��g��?~��}��O)�ϾC�b��,��[�&����$�tO �p�ͬ��4��]��z���6����m�n���E��nY&�*D�"��k4�������Cg�j��Ju� ��m�8���[��J�=|9��t1=�����1F,9���1�m?q+ �.#1?R�]jN6g{��i��%�K���p�0�3��9�G�LR����gh(}Y!Y��M*����(�EN�;�@�hY+aT�����3^�	sGo�Bww[�d������GS��`\e���������iV;UP'�b����6�l&���л����6���: �h��k��G/�8So� �{ ��|�W�������
wX�(7��g�k(J�|x�@��Yb��<;�����=�`�!�=Q�?�sw�nT�����痣M�=���Η.��fi�'.}m*~���>W% �J!��~�p�d{}S4�6Ɏ6���b~�^ђr�S3N
Ǝ��uo�)��!b����l':mG�1ޫ�m�D��?�5���W�<jŶ52��"����Ց	��/��T���l�i��Y[�C�����{E��%��(��/�&��u>�I�>H(\�b����Ӆ�ڑ��{f~(����K�D�Z]�"��m��}��o�ſc��,^�9���eW�' �Z���v
��Vά�N��BrU+ry���⨙VvL�tB��#Ƈ��|t���`�	K�P��GDE�-����-�Nsp���%Y��s�C%K�����6�PF����@\���P��}?��gb��-k�c�u����`*��4�rp���6�sF=q����n����m��j�#n*�[�����davY�	��Ҕ3�1��N��ܘ���@qov䀦����.u�	;D ��ٙ���y>���� �M���������{ġ�؊i�#�5K��� �Bu� 5Ke���s��!.�2l��k�50%�ߵ}@˅�R����e�x8����w���D�4�|�S�Ds����vɤ?�Ч.10-�1�z6Ժ]2^�D���7M}q�[&
���O���0�:Mߖ�����%���nl�4XlDVi;Z?����q;.]��fՑ ����L�ZP�}%"e*�= �jZg}$"%��u&N�>}�f�L��OR�1ݗ�;ͣ.cp��Y[k�0�_p��+�ZȲ��a1���N&�&��x�V��ȟ��DKP��䤂(�in��`C�|�N~]����Y�<���!�Y��}x��f5Fڧ�qu�X<�?G����w��C�'��g���מ�sՑ��p$	�Ĺw��|��L��x�1g䝏�T7;耚DA��VTd���!ݟ��(�2�����N)0����`X�D�%�/ț�8��0#�EoZ��` @�̠��+��G�a�������g�"�i�I��o"�85X�A�azp۝� #���Q�V��*��^D�V{]�(�r_���w��f܁K��G�o7����;��ֽ�zo�}�"����{x����zk��k��Y�K�C%���03���Q��6�T܎��L&��¶HD�����R��!5_�kԦk���l��>7康�|\�,�-�V)��d߂����޳Q��=e�RJgKYƅu�Y[�����ٴ�1+��|�D:�]��H���%�����O_��ߺ0յ��n���W���%��ˢ�]���W��K8��ۏ���lE�;(�\46Q�]M���h�f�	ӈ�leL���5�bj����j� y�-3�Z�\�V�=� _�n�OM��]�[ E/�#��9���m��̘e�Z̺�Bq
�%�U��8�'�K����9�T��i��)M��@��+�DGaI�[!SL�y������w���6�׬�nE.�0�w��%�t�ۚo����\�q���[���#(r7CfI��܂�Suބ�NlV�`����W����V��y	��z,��� �;D\WQ� ZXE�N���h�Z����e�����m��k��vO�Ʌ{���_R�Q�5���U�$cg4��,���~`�p<�Lv��5�)m����/�O�Kդ������Ӳ����L�Ռ�S����@�8ƷuӸ:ԑ�%�M�Xh�.�2\<I�q�l7���eĉ
0r;�C���\s���[_��U�b�x��Dn[T���GTMz��O����[���VГ�)�,�5��(���i�K�Ə�G�Hg<�ˍ��F�Ƴ��˙�-�~ ��&��f�S���l���������#V~o����D{J�h��C׿�X�`�B���mT��F��@>�D���Q���h����S�g�*S��<��.�ֲ]������8�@8sM�@L�����l_����W��{�:Z��&�Z�8�F����J$��m�iC�R�?[�
���.�k
b�k�X�[VF�x���^�U:h�K�3/m㷼-����VEh�7���d�sppnjz��ӛzTƬ#3!G2��!��T+�cJ��e��m�e�ke��p��Ũ)�\k��=KS9ͣ	��0p'F�]T$��k݊8#��΢,mN-��=���[f��7�dt�Y�}hhVDS-�����C޾�f����}�f�D̮9�p��^T���qE�;�S�<�Xwꛬ����<�JF)�<����y���b�o��0G�o���Z����9��[jP%��HwF�A Fˬ�aL�<#,ѫb����ХA�Y������F�!�G�b�\E��r���gT�����T�v����p���'�*1��>g��A�y)�^dI���w��Ȃf��9:��s�ն���S�S�X)�t�'s����8���mG0+�ِ�����?�坈�'��ܶ��I�"�J!"2��� ɭ��et�0+e��d�pɚ`ن��c�4�P)���JuyҰ꯬.8��D���ߦ��'ZA9���TB�x������A���kߙ��O��)	^ꁳÁ� ;!x�!`;ѿQ�6a)��2��:���.��<�iN�
��8�D��!
�{��aV=. %�î�"8�-Z�P$�BD݀�m������2�He��n�1�J��H�H�> �-4-