��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��=�P��q�n'���}6𞆤m��j�I�� ۊ�E0��`� Sگ�v���ҢWs��[3 �z�XW��И n���W��PDo��Fس.<"t�bhS��A�P��M�5�I��mw?�h�s^,�O�L��,� �}?�2���VQ�)��.^tFU��t�{:�Ł��1���t	&F\B������V���\m��cޏ���� P��k��@� �f�g����gc~=���#��/���E�p�´�
9�o�j��B�;;p��޶jYcDp��Uj�=�XR�r��*��i�p�������(#���(�$ܓ���/}	����A�GUś��<�n�����h(��B��,����s&f$A�o������܇b��|#��[��Sk���OiF�����h�8@k*_�5I�*��+�-<u�&[:�:����f���z�X�ʗ�;̑S��O����SHo��[�kW�t{u����\���[J��6����_�jN��.��$%3)�ĨQ�:�n�Y�k	QZll���E	��=6:��[��m:�s^鍊>�Db���~����{:ݦ���|6c��V���߉�ٷ��m"|���W{�`���e.y�E�R�b+Q�F�uj��d!v*%���~�e���<��D���K�?��'�������&�;�:C�]�v����� ��Qۈ�A]�i�ni���$��ިȑW�L�%`�?��=vs �p8��Td/��l@<�K`w2��| �,�kp������K�<+��f	���Lą}b!q��� 0�e�N�g�PF�����2���~[��j���r�MC��]h�3weq�ƐRe����l �Rk������~Ѷ;�0U��"�l�GC�@1��|�r�Hb.hS(����`�dQwn!�~;L˫���߄�X��ďy���8�t\���[v�W�('Ҽ~���'W��~?��^�7S4�L<{w�ѫl��+��C����W�JV�q�=�(*���>Tp������K�iR�;7���6_�	���pE�iܽ.����dy����s���Jb���:���g��!ڿ��R*	�Pͤ~B�@�4�e;����+�Y�x�c�OT\q�:[.�0�3��%�qڨ�A�)����(�9:�PF��D8ƹ������hY��=r�f�Y$
َ��IXt^��"�1Wt�yzӟ�Q;�z����&K�F�%���`K�1�)����LJ�1榀[fz�,@孩@��e��FQw�K�t����6ȑ���qo���]s,���n18�-�J��W��l���m���w�p�_{AX���=f#�iI(4��%�P@s�t�6WY����D���Qө�Ua����A-\�b���&�Ɖn�����7�=�H>"	�#�0��k�>V�g5E��|�b��K�Gk�-�������4�35�t�
�R�p�$ƒ-��|�4���n���S��a��o8	�����אA\�6N���mL�,(L�B�����%G(�a�`��O�}�sOvz%���l��im9��D�m�ߨ�;"���98��܌�:����[*P�VR���@	��,Ng#l�r����v���� ��A�2��E����p�1���щ�
<�C!��I[�!gŢ�q���gf�)<��
�@�tL�����1[	�J�W��W��V�$?pW%oｻT?}�s��y=3���Ђ�٤eYϥ5b(M�ØbT�����#�T����K$L�2?}ǖBE,��k��E�J��`�c�����^g}Դ�H�T��x�"��
D�D�V02惮�4����ª~|c�f7 �Han�#Y��WK��h�X�9�s��z��W6M:��b�]��r�A�ļݺ�y���>���>㓀ygr��b0[c��N4������F_0�l���[�ux�D��z����3��[�-���c��F)�O�H�,
����?�Q�.�ZQ���w'�%LA0鳆�Kb��u�	�?��ƨÍ��
��;��M��\����T��/������1�K�ķ`��~��a���)Dk���͜R*�ZQ��c�r?����KS��>��3!�ȌW�Q������-�z��"���u|��1�{J������4e��_��M<���f8x%۵��a	�Ħ��Y����UTn�ߚ�jP�ag5?o��d� ��f�Hf�ȍ����E��+���)�
����>����}���
�#� ��8�m���l�4�[1�tb��'Ow��x��� yy]��/?ج2�T'9v�R^ȴ�𙘓���|�вwu�)[����h2�|������$�
T��<���騆�Pq䙦tr���V�*���̜�RY�Oj������;��n�/~���4�AH��lI�����$G�GT �5O '�7�Y�e�u�6ϯ43{���uշ�"�+6x,��
p��<�E���oݽ����L3���v;Hc<�B�-C���G 6�<PN	=���JG���gC5s�Q��,<���/���a&���#i�Ĺ�'�R��J͈S��	�N��~�SC���E�!`�@���~kO��z���r�%�#�D��1Ih�u�썧V���D����xJ*dn��U�k9��~���!���}fW�WR�B3��"d'D�=M|7��F��
�m�O�ԝ7���9-M���l��"�^�B�vX$�`zo�4���27���yf�+^oc#i��R����>�l���&���k5�Tu��dR��C��>3%�Ҧ{��<)��G�����VP��ԩB�s��5�3c,wp��[&+E��������HJ�4��ydиw��e���������S���kH�р��ֳ��7�����-{>�OK�7�������+e�9��|�ӽm�*�����Z �C/4�����@r��`1�:��|Ro�F�-, ��\&����-�6t�L l7 UU�"P�x�1��MP�d��)/C-�r�*��/� �s��u�O&�v�jJUŏr;�&\|̓�4�e}-O����5\��r;x�N<��'܍��.����3&��G<���8��}�s�}f�>�^Zݜ�����a-='?�t(PJrM�|�u�tG�:W��O�eEY���S�4�_� �ǚh�ļ[f�Q���-ppV;�I�佔~5JPp"��/E~��$C��;�X>Ỳ�(���?�t���Y�hQ~^�%��6tkw��־���5 C>G�h5[�AF�iM+�):z���#�-t� V�35R�C�7��;@��b^�F#����EdE'ng��SD_4�g���O�_�snY��x�<p7�lV/s&d �Ԯs��FU��T��U�#�	��}��K`ʨ�{��m5���?�ԑ��g��b���61>����Y�J���u���kv^ ���	Ź{�=��Nc��������.��d��'1/e�xw�s5+?0����t�x�*O������q�7%��Wr���d8�Lte�T�L�,��L���J7��}o9m�J�P���r��rmn���7�?<9��X�RĕP�F2��4.��Ge��IkÇ ���'uGeC�$�����AN�"lw���X��?/�0��w�fzG_#��_�
�[����H{x*K@�ĒH�1P��ϱ6�:�PSt��G�eܕ"�%�3����J�E��j�y4�����ɡ�@.;�F���uX`R����E;���T9��.*��*5�n�kӓ���S�=j)��A�`�j5׶����]k#�i�0/�
8����eG��oȭN�%J<��
�)�GO��밒x�FC��"E~��gm"�VVw�k1��pK�
�=����%X����ܱ���o�h�d���)o��#k/��ـ��K<�C��N�:�K��?8H���J�}���p_"����~Rpġ��6�����"հ�W�Jm��C������i�D����X���ey����bB�Y����w�"մ��B��Bq������������t�ɻ	3�y��kZ2tj�:b�㑢X������,%��qjy�6jx���-	������R��S�GE�wՊ��ds��뱲�3B��]l��d\S����X���;ȝ'O9�t�pݱ1Ƙ(G�}�5w��Jf�`׀�XW�.������7���NLt�O$���]��+��c���nzF���[𿥨Z��Y�M{}ƞ����>����r	Ħ���XZ1O�c�V���a�O6�����*ms���΢Ȕ]����N�:a�J�N��iRڊ~ҥ��\�������SG�JX����OC�F1]b`[�t��:�f����^-j�����S�b�e6���l�!�E�}S�	��>j�U��&]E���L2����q��aI�����u
�L��_���t���o���d
���B܄˓�L��g A����������Èb[U����P�z;�y(��Rj)g�ʇ�Ou�{_��������D!�`.��C?��6����I�l$�����V<�9�+u�&nj=��<c�ް�m ��ő�mID
���%
�T{M6]x�V�m�o�qPV��p�����0�8G�}H�#m��se�e�?=��U$��w�N
b.�#�TP���~�n����a ���Yv��cJp.��:lFS4u�C		��z�Sb5��:�us�?eKk{ �h�c��H�"�oJ׿Q2v��o���D�B�g<��b�����C�eR?CU-T��2��}�cP9�!C])".�_�z����L,VE�:�]�ڢ�H�����	R�q�ꀢ���#"(�m��q�X�*������#�?���#���y�pW�4��<RU嘾(	}���L
]�ADG�:mKd.ՙ���vG���c�:�������{�8���M� NzT�W��TvԠ�{`J�]��&�E�c8�K�T΃��z���:�*��!e?���Sw��0�I����z��~��ଂ��!#�. X�x����A.j��!��e�kEoi$���J�ѕ��%�Yډ���R��~�`|�}U �����dʶ}P���O,��˙�;�o��5�Izi�WL��mi��\A7���q�˕�7-�20d� ��������U�q�!K!,�.�_�G+�`�4�C�o���[�
�s��iosx~3F�ϼ|9�F����sG��T�g��0��R]�����}��;�̭{e?,��>�O��O�����zNK�
�]h�X����?[ْ!߼ğȆ��X�ˡ����>�����B(ŜN�n)5�DQ�?>�������HdZ���+�)�TbK�$�=k�G-Z�t
_2;���%�U���ˇ�sY�͊��0�!Pp��,n� 6&��F�j�'a� �0F�s����:� h���&��&yt�[q\�	'��J�&�/�?H��Ǌ�I�u�Pו�7M41�%G�`���0ҋD/M����.�	v2�$�I���l߿�)FiS�ҳ��/w�"e�i[)Z��P��Qy9�l�n���7�p;G?P Hd� �
��SOf���<[#0a�Ԏ-��P��O^L�K���a���P���z����x��:#�Ú�J3�$��I��lS��\	#��ɇ@��fo�,&א�p*��VJwcDT&�o����0v�?\�y�R�����������vEx���%�>g�G�	�B4�4_��.�巽�
���`[������4"�ʢT�t/�&�c����]�Y]�2����9�`ZQH�v��L<T�"3v�+i7��p܊��� \Pa%&h��։=߅�e*߽�	�%������_���;���4�%�B������f� ;���q[N��؃ <��`���ϑ�lJW鐪$�}8��Lz�O*y*!��E�۞�^���-��1~Ju5�/�1"SІ!������3Յ�{�v��;�nJ�I�Z~�*%����*��	�0�+���d�TY����/Nl�|��lA�y藣��J+d8���ٗ�� ��<�p���AK��N��ڜ)��J����N� ��P�L}����Χh{Jx4jDJ]����y������n@�xd~>��T@��J]r� HQX��֩b��j~�&��q��>�I�DD�g y��>��P��dx�������<4#�~��n���\t�r;n�r1��g��#��b�io��o��*vHy�#���+m��|E9�XVK��ִ�B��ҡ(�#z�o6��,��h̪�2�mc�5���א
C����.>p{��Jd<C��5�H��&�(x�^�q�~Z��x�)�E�� K�܃�Ǯ罆��22��#l�z�k��YT�*�)�n����h��%?Ω��GlO�$�U a��	�[(КNF�LY�.q%��Cޠ���3ވ�B� HzY�x� �BE�m�ѠO6[ nًUQ�zR��I� ��IX 2i�+m��g=��x�I%�nר��|��ڊ�+e���>�8J�j�ܝ�6.D��0U.X����T`ri�O�}�9<��2�A�m=c޾�A۱ى���wT6*v��-�@(�#NU��"Vp���(�o���ٓGn�����CK�/�(���[�es�K�l�X�:�I�E����an��ڙ��M�@���:��v5�a2R/)xf�!}ʓ;�6e�atKJ�wg�*%�q�����a��F"ԑ�$��Y�@����k�+5ՠ����U"�c�[Y72����X|EGR�ؤ'h�g~u�4[�w��w�Wqn��u;���ю�#ׯ��x[_r�q�?5K�(�0ʱb�ɲ���X�΋�Ck��_�<��d^��-�آ�!�Lj�2�EOV��Ǟ n69\�k�]',�I��kc�L�H�iH"(�7����D#��Q�u`YKJG"����	0
�Kf��{;�w	�RAy��I(&�!����rįxf��2F���*�NX�����O�6']�s[(�����r��<�;�*I�IC�:Y"e������/˹n>0ZǇ��	O���>'�"X�Le�� ����a�/��J���	�i����[�]<Q6�8%������=��^��b��Q�f&�I���9��ScKUz��}�Y�v4�@���a��{Xlz"K���������d�D���<�vMAˏ#�o�
N�?�Y�0/�����ٰ! ��������aX.�?�r
H��T=?(%���ܾ%���c*�>����HƸ]{��lC���t	ۋcz��B ���Z$Nb�תxoڃK��f����ߋ#�ˎ�{�ˀP���|��0����9��秎��ҧ�����,⥰�"�������e'�^I�my7w
݌U�Y��ER�
#�ž�_�Y'ljEC�_n���B�Sy�r��X��O����[��x�F�c�/x���w�M;s��k4_���%�zjg��U5�2��#$��i �y���=���89<����}'^+�����0m��V9�]��j�B6���8x��0�sxN�<_��f����=���[��~���'~���p=?�'SM��E�}��X���~�:1��ɜ�}o���H'+�:FK࣢o��*�LG�I�n��	����S�AZ-�qػ�ʼ��
�,`
�O_��@"t����=�Efֲ�ӄ�'���U(Y�n�e��f2^��A�)�T$��/�mA_x� 	S퇏����}/���S\�m���y����3P����@����M�"�0�|���X�s#�~S3����J���U�{z9W�iw�-��v����lvS���P�!��%��C�&2�o|rD,�er��bN	Ʊ�Q�9�����Ҙψ'�审{ӻS�u[Aԣ�x��̴#�.T�؀�([w"ݞ�m�D��ڱ?G��۬iY��l���<��˨�o�C�}EWkݝ�ғ�%����<��#wq�|zǘл�b�ݨk�,0�����^�%j�C��������9�#��*K�=��Z�#�<%(��>-��v��/2�GG�ԥ�F�\]'�B�ׁ(�juj�њԊl�{�`}�
�b$�{�Z��Z��{�+�_X���|��+������|V��Ha��K= jx��	�^ʤ�<5	��}I��[z�>]~#��N~��-K&��.������d��#�� 44�DZ���q��ˁ]8�vVS���wl�P��[r��S��rQe�"�A��?jU>q#��7����E�w��n��9�:o%5�(̸��EX3k���*�0���	����b
Emx����0{�@����l��h[�ښR��ovR��"Q���#(Q�W�%.��!��4��I��S��j�5�K��[��M�U7���׈/�7���S��Ԑ��o@��7C��?�@i�	M�4֏���4e�1�)�EQ��)�o�5Y��0� q�S#I9D$�ҦI�U:� q����lƚ 1T~�M�i�}ڢ�1��A:�ؚ�ak3��w&��+�����-Z������i#߸���Z���r볘��fW����U8EL��m0�ض&d;��]��E埞�-�����̶[$���8�ϥ?���g�wy�tP	��/W+k���D-Q��iyg?������r�?���9q���D����Mc�
a�7e�=E#~���g4�:4�H�GEC�u�/��>dFxy5�s�8�J��@-I�����t�[�͟oS���Q)�do�q�Y�����rn�^�<a�xc��W��0�T�9��Y��+b6�q��Y�h�`ap�:ʲ�����WC��I��B�N�� ��{tü�]��I����n�N��Н\ڲ'�J���T[g��u�0�i�7���q��L�;�i�;�~�p.��093=�qg��;R���rM��W۵�[��Ň.�Օ!eQ|�5�'�zLbP�{w
�����mXbC6X�e^���f"X+���x�-�)I��h�p�g�|��������K��.;){����d���7����u�����8:)��y	=���2/S�D������Z�PaT�~@�.������{gw�mY��z;l}Ud��d?N
w��^�r$�5�С9�����p@��E��\�����q����ua�'�[r�5pe��hJ�"��t^5�h��?�&K���wM F0�m�4����3�&����V����}<m�-�NzG�������&�<Hn/��M~�7mv���a:�/q����ΌG�3>q����i��f&s	b�y���pV��,W� �$�jw���+��8�㽞.�3��ƅb�;tN���0̝��샧B�~E�e�����imć7'Ϙ��|Y�X,"rOtN�䫧/��e���m�94q�����W�݋�q-��v���^
�D�}��6���C�'_r_CYR�-�2��]�PcC�?��,@OKSzG7ĳ�כ�2�@�󋈑�[K�3΄�:L��wT��-Aw����;$2�}-aϨ6pʁl��mip��rlLzNڮ��6Z:�EQ�1�v��P9w�'���X�vӇH֗t���w^��� ^��Z�id����)b�@L�����NN������@pJԭa�̖��y��?S�mT`}��w�@��Uu�a���c���PG��y
�`����~ ��F���x� U|�C���?k��>�������8�N �a��"�^`I��v	?(��`�k���ez��4ӥ�&$�`.��K�0���<���w�s�/��by���,�#��0XW�� QTy��{\���N�*8@Rނ��ܘY�0��a��@�qA�~�C�q����K���f���1�w�L��3�6H��m���;kx������=Έ���:����7{L����a�`��V�*�!րzMg��L��W�FyT����\ 
J6R�����_�'5�9��*����>�ܻ#�J5u�V㐄���DP�
�Uv�*0b�En9)��ٿxx��#�d( 'R�  %eC�Ef�,abҡ�:��K'x4�̿��t�F;=�o���rHύ阄����t%���{��%R+�P�SS.5�����phָ���\�}C���7�[���P�("Lq]W1Am�	[�I���<��(�]j���om7Uz����al����]�&A=�8ח����R	�x-��{ăQo�"�$lB�<�k����y!���[�L�k(�˲CN�Ф��X��7Q�ʀ��  ��H�G������WY�e8���B�ǌZ+u�U�*.��M�#����*������2Mi�B�vĩN�H���ƻ���QQ�9�b�2'��K��r������mSW}���)F�P�%<��p���Ҡ�C�^}!l�<�!�,-\
���Ի����$�+�)��c��_>��,���1�%Y�M�y^i	�On2^�lGj7R��-��b�f�L��Z<�9��. <���{��ג�cH��*U�t�}�{B���8G��D�n�`2sx�^�j��u��;�`�r�`O�P]c��
^�V���Ď e_�K�rN�WZ��E�Dmy�[t���e�-0N��ꙇ�0fK-B�>�n��!��RUr]��Kṵ%B��wH�4�(#�|��l���Gs�y���`���đ�|#��z�����r؊�{�ذff%��r;�n2u�#} ���
����G�h��>���A���- d�ZU7K^�^�-J��2:�,N$��)!���� ��R�[��ۡ�ʓI3 Dqz����0�Et�	�G[�z�<d2��'+g��5�~�i$���uX�q���/��0�
8�������m9M�f�f��l]D�EG�ZuTv��Ty�E.�� �Cf[B�ךJB��Cd���ឳ��@Le�Zg4�>����u��o)d|9��'�����I'�z�6C�����両Ro,�ʣg�?����Og1�Y���!�ĩ��m�M���4
A�]S�K�Y��b:�X� �)�d�
L���+����V?�u�!�1��n>V���o2�S�ڐ��O�N�E�&���M�͔7W�Z��8Ekqd�O^�U�_޼f�b'���>7����Q�lJ�k��%�{a�8�N��n�&�}#C;��~#!ka�n��5�G���h����6�6@A�~#�Y|MP�J�s�������\)o�$�M�s|�����(J���f�I=��NJ��u�hCI�??l��^�
ba^~��,"����%��|a�=�����'��\��	�f��A�?�Q5�柷+0wpT,ƛ��J"S��f3�r��q4	�k4'�k�W�4Y���FY��'FF#�#����7Rzoe8-Z��a�c��l_ߙ��}���J�r���lel6~G4^��NtR�"ܢ�P4�]���[����x�:o��3n}�C��-�>��X�]
���x4p�t䳢IcFK��nk����-g��xz���3�,��q�
����z�h�T���"�Z
��ZU����֌Z�����Q�����-�}�a-�R����%Y���J�f���`�P݉2�#Ne�`�� ���թ��6���K��\I�(ހ�c���h��4p�Bu����MI�ڊk|�O[�ۅBO0��%:	�@�Ss�E�[f��zt�}R-g�2�����}(�s�[���7޷F�è�����	����ʨ}�u�+�eKQ�8���I׿�=F��IEO�-�?�ė
���e�(�7�`�1$�]+���W� е��rJǛrX鸪���x��Я�N�nG��f�����"�|���N{��4��:��5uFk�6�H�;ʳs/��ozG&�II$��bt�@_K��DwY�y��f{�Eu��
&�#�yК���iBTVD,�����o�y��V��7�e�>K�Bc~��+t-;��"t����#�1�c��l�(��X���G�DSVd+0}|��C�~�����a����[8D��]\
w"�,#Rx���z�g�
i�E�q���Im�I�����
���>����70Y��*��4O�(�sp��%)���O�ٍe�CHPƦ�J��ˁ�i�;�x��0ЛTΘ��h���o�ۜ�'�z�U��$�X|�Z_�h�{�51����@w2��W�bi�x��Я��q��x#,���#d�e$�$��05?ͅ���;lU��>��%@S��S�W�]�?`�]ܟ� 67]�~�,u�y�}A�h>N;l<�Βtc�8O��
�Y�������4�VPN��7��J��J@K�kb#-�p<�<�gx~+��K7��\R�AU���{���,��^�����鳆ض���#�o
b�@#8�� ���n�����ہ��Y䢎<���$K�Oت�4��]�v*��흍$���,BS�%��X�i�i���%��� ���k�p����&��NObP씜�p�lZ]��zGq�C���7y�QP�� ���0�8�і����l�O2���D��y��n�L�`��}ϟi2z"]>��!O��A�F���t�^�����v��e���0��Ȟ�_�_e7���ȩ��&Ɋ`_�U�%���Q���rrq�骲��:�+p��f������8�.&�bd�g�a`��Ĥ	V�{��/��
0��u�;�=bA4$�"LH[�1)���wYQ3��*<��k���g�<!��~=<�f��7#!/���᪲���|m�v��{ �N@��܊�w�g�ɵ� QVl�Zݬ}�P����i���XX>W�z5�B�r������N�]��b��^s���i���ޛ~�q=n��B�ty�����{���X��TH��P<� n;��.�G�y;�;��;l\�!�a˗iD�V���i�}xF4�ܞhXoD?�<���c� -!�)|Y�8S���VRa���&���f�/���y�*�y	�QS��W�|;�t��� �F�l7+�v9%M�*���[��O��|�jsxl\���g�	:G�/���0��ѐ�+�Uf��U]�	I�g���ste�Z<]^R�I�H���e#��N��1�X��H��ѿ��A�pU��{s�����,�=;��`s�o�Ԁ���	�@��.���Vvl[�ɰ
?8I�I1��'�븩���_��1eh��4ۂ�]\�s�cD���?�'�Yўb�3�?B)��������^\H��j���DT1��M��oFa��a�����V�P�"�qD
��k+�6G�g ��p���9��ܸ^}�c/�'�f����L9�D��fo��2<Vj�u--63!9	�:~�.T����'}U(����t~>�Z`<	��P2�������b�ʨ bD)#�Qd~��8� ���	��(
�jf�B�@�g���m�Pp�����I�������FX�˯c��	IC�$���s2�S�1����˵!\���z�º?,!Ǽ�̧�_��7�qT2^*+Û���:p?%��� %5��oP��Mڒ>>4AL#lՏ��Dt�Hٽ4�#9�^� ���F���e���B�:�&�x��	�
�D�g[��o 	d��^-܀��0�Q���iYX���	]��.�.��yR��~J�j`��b�%��Y�,K�\�ۿ6(�@b���[�R �����$���xˀU�r+u�|�3�K������_���հ&�@71~4
q�Qi�dŽpG�F����ֱ��(t�~7�e���Q,[ST��ɤ0���@������C��!� (
8��?� bF���^��RW]�����X��V���=��٥�����w`��z��Z.�FH��g�o�U�^5�Z����5kl���oB��ةJ%7���N'/�Rr���y5��o�G�����>O�X��l��Ȳ�����u�hMвJ�z0�'2�9���W��3�p�'
���CZ������3�3�֩-d�g�-�6��Æla��^fy
��s}����+���m�a����|���u\��qٷ�
�Lό��)���^/&�!W�ۜ5{1ǐiX��r��w���&@b�����U-8-�f)*t�ï�"�g��U����s���C'׮O��H�L�P_l:�Y2�6͏��i������Hs��\h�+��C�n�9dY8.���'27��@ ��)���c5�kq�d��U�٦Dk�����(�+�b�����W;3�#DϺ�4����OV-����tT��(�?�_�6�<����Z`�(�Z��./�X�"]�
�@�H��}Z.���lW	��N�5w">���Y����	N�s�Kl%Ԇ�P'� �b��2��a�Z>����軧0N��)_�mY�E�%?=�{���H�Z$��V�YTi��aH��0k��k�%0V)*���Wucz��JSV'�((m��_��ԯ�`fPo"��O��vB������HP���x��w����;�bt�l�<�����/Ѝb��\-ԓ��qk��
D��e�n���x-H�l�v&Z� I�LVGKq���5c2f��PU1���a�� �f�	�撢5��k�ʋ�E��j��P	}�F�ɟ��o.Fe�<݅36�z��ۺ��B�W���
�%g;kt�r��ﳗC~�M���)����n��M�Tn��c�[5A=HA�Ӕ�����Ӎǻ9�B:�� �t��ə���{���/#�w]_���f�ۡ�����*�+�#��~;�brB��YL7aM6\B���rrKN"���2���H�ʬ�j�*���G���Ҭ>��<��!'M����{��:�d.�y6&Ļ��֊N����1ؖE�Kb4��4����|���i&�53�@�l�\d"ޕ��L�- 0ص6;����d��A��8{Ռ�l3�	���c/u}H�[ K�k�FǸ�Q�B���g�\�7����I���8�����H'b��%[�R����u�Vfn�@^B՞�"��>��٦����Ej }x���{�$��:��A6��8�1Zo�D�U�����;�mIz!�R��.�w��f	���u�iڻt����K*9��p�n� d2|#���g�>������q��-�=��������2�"9l<8b�o�a��=ZĤ`��>R��ե�<�U�a�"�� �]B��G��C�լj��GϚ*4�Q&��Ix2`�b&43)��)8~����t�*N��8Y��"��[�+u:́K�_䦷�<\��)	Ӓ.�ǟ|K.�����o��2r��+�k��'�A�D��o¾m6�8s��V
)�-�J���PͲ���D1,���h����o[q�����)���03)�Pt���10�V�C���o�Z`��_�q�fU��������/s���,ˆQ�Q��xa�ƕh�،��w��1*L�@d4�zB�D�bm���x�j�l9�?����	]2��ܚ�w
4���L�"��M7*0뗍�~����QGC��7=���+7��r�ۨ�ȷݞ�!2�Dtm�N�\��ٗ3nc5�w��C��R���G��`��(�-?W�l�\F���E��)�~
2���1�jՉ����o������N�1<�Ӡ�e�u����$'�ZKGC?L{:�4�b�|�k@����,!
�uĖy떍�ޣ><��c���[aݳ�R�7P楶܍��ٮ��T\�M�Y|�ǚ����[4��͑��2��l˺V���8.W,+��4���/&R]x�ҙ2jH�ւ�AE��!�a��md8'��)x��zO���B�r�KR�](�m�phO����#��Ux�!\�m�Y��7�N
�ޔC��"~���@������,�����dq[�ؾ؍ԯ��!7���߹q ]������o����֨�������ES}l�&U��+yL�7��[g��s��im}yS��:��f��3!\��Y~BCU]>T�Uo���1$iz���:���7�CD4>�T�x{]U်��P��i��XG��UJ����GWU�Go����P@e�XCZ~�e��S]�������O֗���$��Oûޟ�a@�5����b���*�
z���0���2P�<*I��e�����շPngyEX�-�7 ���[���a�=�q��jpk�*K�U�s���S�.�NY����w�m(�$-�e"����?>��ei"AS�\��e�%��E��=(��z�7G��v�en����l�����81�(�ʮj��9����N�
��1U�\l<j)F�N�u�����FmteO4]s?J�n�' ���q��
e�R�מ�=�:�Dׇc����1���}{m��hت\S��p���3Wx�;���<���[�ӍS�?{]�,��&i���Fwi�ȍ�p�u�0I����B����=�s[avy�4����N}�|����_J3�ch_��OP�uF_�	��
���ߞ8�Ұ�=&�mj�Txj�Q��~]+E�2��V�i��Ô��5/A��|*�=5$i�؅�p&T�h9.	{q�N�~���?=�8 ,+p��"F��9eܜ�Sd�Hv�����I�o�,�ۺ���h^�8x�靆p��`Ҡ]�%��O8�B��YmG�l�@S���_�_JJxBl�H�d|�v�ُ�{�F	mM,,a�����`'P����|P�2�������p������x	��q ~%z`��Rk|�k�S�M���WBx�$�z*ί-F��Q`��A:���bM�0_鎢]U�}y;�?8���ɟ���P�f��&~��.V>.�nt1���o�QE�R�a�Lwk��3Vz5�x�U=.���@�N�%��m2Q�(T��R@V	�!�K
��s��5u���&�S��K>G�ܽ�ٵ!~��bo�[TY�M��RU�Zz���>�,
��D�;'�͍|�ͣ�<9�O7�QI�Ɵ:�W��.͎\��|#w94��b���hg.�DN"�o�]!�whT��C���h�]"`=�£P���b|Bv��j`˺2�����e��8}�����龜D_�y�"���wX���{�צ�LV"X�G`{��׶`o��z��Z޷����� �0��7���`S��ŀ�H�#�Nn���jˤQ3����y`d���P����rOh�����&��t�[I���R{a>�,%
�|�!Q�Y�Ds��� ��5w�
�F��Z��e7�x�X|����*s�/6�U�H2�=���	KSu�� ��J����˔ڇ5�vSc�fo��{��.+/�-�Nr%Qe���cŉb��3=�'�QT}]������%h�*3���0iugX��__7��I�h4�ލ��g���n�	����E`��x�������>PP�Y[TlB��3W��]l��IO�2�[�P�0������毅��b&�dB�U�CHuwR�4��jҹ���g)��>��vT��j��� �Dd����c�p�,�&9�{J�I~��V������S�b ��,"f���!��!�k|�7�ڎ���>B��*�[M�<S�*�R]��M[�)���1!R�-�o�e��H,�%pq:�+_a��A�)��t߮���͚���()�u�6���/	�F^#���2 ��',���q�J+�1�/pQG�#kf&��D��bnp-!��ʬ׳q7e������#�,l���$���a?��.a��1��L�7�<���.�yx0�&c�X��\C�ܬ��>۟>2�v�������O��5��w�K`l3��1�
��3W�%Lp�	����VҠ�����g����ʠ��g����A����_eq/�G?�0�:��G�8���@\�u%��6��i��Xu�	8���oE80�;̣�34�?��=�o�N��KU��H�����)8��v��I\����%�NfTX��G�/A��t �ɪ9Lv����I��T]�+
(���L���l-�o�����i�����������S�kF������y�n��T|>�\�������9C���������,��-L�򌷰�^������R�t�V��|�*wX�S]��JW����NӦ��F�+������E;�$�/|~�"؜�L���(;�i/�6�������4 {�N-6w*�#JK-�t{85�LB��p����!�l��FA?���t�uJ�[(�/�8�~2��ڵ�v<�l狭��+����X 1n�N�`r��mm��2�=B�`V�I��pK�U�%��9���W������C�����ZE���c��j�y� YOWL�ٹT��k�5�r�T�9�&ԓ$w@������)Z��
&}����Q��Ř(`��s��z�-�WD�ɋJ��6��8�a�ʧ�����m`g�G�rW�/�ah��Ĭf�AN�S���E�\�)�Н��F��������*cd�A%"�Ww�Pcw���XԄ0����}���v��Ha��t⏖�W�ߎ�i:3��D���Lk�5��Q�c�9�OruU��ؔ�V�YF9'aљ�7����A0Ş��-\I���ξ��oZ����+-��MR����e�0�IW�pٱdI�W�͈B9�]�ZC��Ơ�/�4BN�5��]3�����I��*��CK\-_Mh�Uvu"�!�bZ�#������Ԑ6�d��&?��äs�(�~� hm�|#��S/��?N�)�Xy����D�bĐ��%��6���K3���9e��Ӄ��%.0�J�>��q��G�a��x���q)��J�����h���"X���ˢ,DY�3�6��Wz/l���=��_�����������N`U������t����d@�����J)�9`�zK��7�����,�qg��2�����i:�<�A�9��q6�=o^�
e2��BU� �&g��;�}��9#+h��̌}j?�C�&�[#:�ܗr4�����J��i�pnc�'���i���9-�g�������7d��R)껣̌���.���p�o�9�݉��i�'ۭQ��:؀�>W#�a<\0��L>	�Ԫ^�-����q�~Ep8��l�3��b�C���JdWA�['b&¹�<OԞ����!�����7��jW5{�?��g�+��@�������G�p��g7_*���3��/�b|ޤ�؀�`�3�Q�bo�p��!!LԷS�3O��.�9��x����-��Ж��s
Β8�3����b��@�PWhFہ���ɝ���;�de@������V�;\�۶c�Ė� 1�f~�6*̐�X���Z
о�:�uc�_ܮgH������6�X�������=��e[������(6�LhULya���������R�����}��l��K���ƅ��8c��"�n����i <[�pqq-K�4��0.�r;3�>�QEq:��/י�� �Oth�&"0�_�e�'�I��	J���&��u��۴��Ea��T��Nv��Y�n�&�υR/��if�ى�}Y��&	 Gl0;B>\ݸ+V�m�r�r7��Z��ż�Y�ߑ
8~1����y(w�0Hv�*�$�ɚ����c�c����y�;:T��2�8��#6n=MK�YYn�kW0���=H\�-\�Z�ղ�G ��pw���ax�V�վul�eS#*C��k�w��h�$��g�g�y&0����D�Z%��H=����瑱��A��cy��dm����5#I�?^FD���؀���g��!մQG����I���b{�r�3;�<0*<�r�p�	yB�D:��^�*�fܩk�}��U���h��U�A0��Au*�0�����x����x�?��/���H��)�l?��l}
d��:j���b�=�Z���)?���Ȏ�֐kG!���Aڃ۩����F�C��f�����FDF(��*�H8���ɟM�o`9m��ǜ�i�J���v	�ۈ��4�,b�&/�>g9��܊��ob+�+����0���I�\iOvz�4�mZ���lLx=-�_��P?zXpd'�/C���iO�"ye���ۦ҇�cqrmiw�+�[/,��+�����E/�/��)�q�9%F���X�;��i[|J7q.��
��+z��iy�ّ�j��U�.��A�FT��%m�QI��uw�CH�D�}�Jϡ�`֎��P5��QB�0QF�
��\�A�S�&k���-ȑ�;�Ѓt��W��	���W��X���/-��{�~�y�y�٭P;=��x�[����6��mo7�|� ؈Ο^�z �� wb!p|����;���e)��nG��9d8XV���maϑ0t;���a2ʩ����������0���Hx}�m��H�*�V,�[TH�]^x��LK��+lë��Tۡs��(<�.|Wff�9� j�阣B�� x�
V��S��V�¡���R����U�`��7��n�U��Y��"�G<��R�s�{-����x��?B�#�#�V{C ��H����B�C�퉨�C�.��Q�Y����Q�ȣ�k\��j����#�YS�$���Aʫz��")}΀	���'G��&�c�
�ȋԒKO��p������w���ň��L�c�7�ΙR�w[s�� ����v���Q{��\���u���	 G-=�;���Dn'JC��/���آ��.l��%�
`��TPX�Y�Jz�S���I=R"L��L 2<k�V�=C�Q�6�:v�c��GK�E���|g<aU{k��^Q�C ��:�\3����r*�!�Hʐ���������:�̷��D��3�-,�JS�F}/�ÙLl����0'�xc�Ϸ��{,��
h���Ϸ}S�s��Crc8_�sl)I�m����#mo;�#W�қ��/���ФwiDt@MGm�xJyVa��
�Ϲ��0�n<�<Y�ŭ�.&�xaY�B�LAdFx�n�����A̡g�r/�n���+��;g/�r-���]t�|d���'{ �b�&Pe�w⁩Fq�r�B��m��s��&�=e܊Ԫ�zs���~�+�Q��U�l�U�+�.uJB���ɰb�2z!$(;�G��\/��'I��ao?�k7i�d{��ew�qr�J]>����ʵ�MV�̉���=;�%����[�%�|�/� |�	|�)2��@[H:�"�=��8�u���:I@M[�R�t��)� J��̵����D�Q
�������~�M6�1����,����T��ۃ�,�(Z�X�d���-0���R�(ټz�ڿS
���I���N_ ��h����W�
�i�[�:P��Gu}���ª�]��q:�*t��W&VBP.�o㼿���|�X�P��x�"�ہGb�~[Z/Np�5S�*ه��J/%*3���xo?�����$tY��)ҶUAxj�>ZX�\!���?��_��lo��߳���8�5@�ā*2n��C%\�K�$��F������*[Ƃ��¤}�_:f��������H�BzIg㬼C���*j�4��6��Kߦ>]rI�b��+AW�K`o��|��x�����+�S:�L�m�ք?��GH|L�V�3m'�Q
��9��,\Z1ړ6K|��X��/7�;ϐ�E����J�^	�,~p���F[�,ӉdkuD'�;��.�|ˎ
[M`���LL��:��Q�g&�{˜;g��n`~D}��Ź'�"�:AA|���Ԉ�pz�l�����h��h>�:�PހW}�������
�3/���_���IQ�j��c�,E�*��֜;���6�h��j�SVކ�L����rk|j��<�8BV�{���נ[������~�#;,&�	�Oםt���c��q�)��w�z<�n[��#V(�$������8Y��!��+/�-ġ������s���S��ķ�F�N4֘�[��d�8m�Z�ͣu��q+� I���}_�_[7?_i���Ԧ]6Y��
*Yh���ʢa�@5��l�?Vն�Ama���/�rz(/ <�6�߈�O��X|ۓ�X�)��i�l�	&ۡ�M(A~*;�n@�>8VƊ.��!�r�^���k�י�;]���'1����՜���R/W�?l��#�P���ȑ��Q�)
���?��0e�f��v�#;�gL�z&�B%
;-�2����j��A����H:ͱ��mbmg���E���i�ndw�B�;|�=��՟�[�f,��s�D���{�Fw8���8�
���ǰ�	e�i���I)��įt�P��>�@~<��Z��a��p_��$4mO��)ydIW����µ��P��97{s�u,�����;)z@�pB��������H����������N��l�*S1>�x��v��Rѽ]���7��9�X��:���v�V%nfث�Y7�%�b�=��Bl�ܙ��ٯs���X��_^U�̮�6�8k�?��G��Ě�;��'���
��&��������C��gL&��<��c���T�5�33�ʐb���=v,�]�u���� ��`x�Se�$z@�֭�B���p�G��:I����A;^Uy�}�)X���tY9^�Z�ڕ+�;oe%&�YhU���a�+I��#(m�:f��~@��k�۽YK^RB�ʺ�`��n}���&4��s���$�9S�F��4��J�H"8�ѩ֛ZW\.l#\!��u|��}W`�%+z1�_��������}mOV6���o���&F�Ϸ�4�Rd�\�~*���$�
���l�%vn�ο׎�����<m�_�a�>N��|�[�d<��<��9k��F����J���{���k��e6!*
��o��(��4{��{���5]jg�k̚W�u#|���s���~A���Kܡk�Ѣ�:L�\K`��O�JG���QI���)>L�Kf��G��/�� �I�>mW�M86P"��ei��8��B�=�F��r(� �+Mռ5�43�)q�0�ʷ҆glt+W��'�FC[?�p?��F��Fu����D}��bT���,IF��=��JT����+l����w}�,Ϯ4�=P�(M''��f�x��zE�?�e���;��[�9蓴��KU� Ή�q���-�K�>�cdA�z�b��9���}@�j��%5����wtY:� KA�{�h�7� �U%����ύD�\�Sڄ 765c	�V@���3\d�ޚ����+)"x�j�<0𳂮�m0x�!*#�2Ki�mL�7N��G@%�y�ŀM��8"�(��}�&5�K�������4��y��yl_�H{T?�9�P8W�|q�W$��XW���-`�#�{�y�����JJ�D�+�g^��0��b��
R�8w���>�I�j���@lU�r&ʍ���r�B���Ce�L?!VՑ{�Z]�ʔ�mQ�����DG]ڢ�6]�D�'��������n�?��D�������2���#�T`��g��Y4��ǰ]s�W����M|��ț8���akjy�s-�⸺[��^2k�ƅ���m�H�hp�A�w��5�؀+hL�IJ�o�P�*�'gXQ[�C���t���'Ao�\��zs I��q�m��9�M����XD��%��}>B�P� aQ/8b
����C�c��pֻO���]�<G����+�o��:�Ս�!7c�E�˴$?Z��p�#�}wc:�b�?�^�G�5�6��WWg l
������=�Vޱ��R826�'Ƈ�&x�&�Q�X��e!l=c)��/�p{4Qq��ڇ;2�/E�L �^�VD�G�&��2Y�v9�����t�-hn��E ��4�yװ�� B�sR��ř�qg��?�[=�p��%��M3�_��;��츔ч��<S����I��lg���?��wQ^��c�}uҷ����l�VJ�/Y�ݮՠB	7�M��ܴ�
�l��B�|�o�pV
g���3TN<ѹķ���?1דx$�H���Oi�A��b,�t|w|m�3��p�K������ҿD~~a����?�A���?t2l9Lzƪj��-jM��?Gm@���{��Ef]�.�!|Ϻx��$���Ǟ��XZ������wCi7�U-��� jX�b�^o�[���եb^�����>����rꩢ48�sR]3�F�il�blx�����@�=�`��1:��U��ڽ�O),�=�%pr/�i��lG�;#5��	/���{��)��a�X�u�W
������׳��wG�����Vkg�◕KƭUi���|��8�Qy�^�I��y.B��ha��j����9�m�ʌ�>���'���Fj
X�!�	)N+�W��M���	�ev�!��
�6eT����O�~�*��.���`��Ԯ[��͵_s�C�*yơ�	ٺ�۲��0ɴ>�g� �JUc�.CS�`</q7��;@�xv��+�����h��um��-��DO�x�T����H��iƓϯ���ؖ�.{��ٮ�*��緿o"��v��>��^�h2$��mҸo�W��w�l6�^�Xxq	�*i�]�DH�KF��v���oͥ�����i{>�1��@7r���@r)I�l�)(/A--�n2X/� ݱ[!&2K�����~o�K�HA8+���ML�+��I����_�u�׿��T%MznF�	�@��5�Ub#'Y
!������s��Bnt�@��,�̺-�B֪�ƾ	e7j3X�hMyc�7�l���?�z�My'*B�C+}�s�6�"{��J��,6ǘ�W�U�$���ji��jj8�3���{<?��a�B�w��?%.P2.��.�<�fhB�5���'�d�oe7�4�p��i�H;�s��r��DSql��u�\�XСP��x����#��c�a`��c�-S��bSO˭z~y����k��Wx4x�0��#^9r9#JzFƐ��.kD�-��_��%�v4��݂e�x\:Q�f$��!�\;Ia�$ϖr	3P�9o��������@��$�FU*��i�P	F�M�/���F�fv�B�\�w<[h{��`!a���\���+���iD��~Q�߸w9(��"�mt�X=��a����IbE�D0O9��S�2EDE��6̌����k(��D|���� �lla"Pb�[�a�VT��'6�e�{u���2=ޓ�' �҄�.�L���(��\�����_ �6�Zl`�����3ju�[r5x�kFѰ��ю�0/�:�E�$"_G�8t~c�
���L���d�m<{<I��:C�{'��&�#c�>��2�J9��)�(�,�<R�r�΢*{�]d[OUtS���L� � Ku���֧$�W�m�X��V���A-CYTJU�k��1b[����<-Hnk:�ìvSL��2.hTpG�+�(}�rj(��f�3�H�p22B�X��I<K�5Jw:�{z��/�k���	!2 ���C ��s�g���$�+��A���{�Fm��Yw�����;��*	@���a�|ns�ڶީ��r��t�ה��r�D) ��
�O�ؼB!A&�P��	�����������&$�6�%����R��N� �8��a@Cأ�$��]В��t͝�3SE���N�d�>@T���8�E�B����;8��k��v��#o߳%����+�S���8=�Ԧ�?f6uB_��s�e�0�_Ƹ%�[�ZX���U�S҂v�qgp������o�Ք�wm�ꔵS�H���?$��o�`Q�p)��ګf<A(/�땨eM�,&t�&N�i��ì��?�JE�A��)�PBc�)�@L{B�Y��}�˙h�H��:�T��T��V�i&� �p@�0`p��#6{�H�ԉy�ܩ��e@}����'��۫�$��{���QD���������rM4HDM\��d���GCs[.�J+:�G��6������+�o_�䩄��g��mV�N�VQ���6o�^�(�.�F�r�r��,q�[����vHvZW�5������� [	Ua4�B5w�:jϮ"��,5	��j�<�(`^3�R=>�HPc�ͱX�<s�;�N�e%�*bV��'Ͷ��&��f�3�˧��,3	s���}���L@�2�RR��_�u`9���y���m*zlߢ��͒�kX�!����@J�f����� �pT�LA�3���|���(�T���j�'���U���M�����>j�JsE����<�k���`]��L�L���#�/tq�����j�{h�x}����Fq���Ja�6� ,�~FkUmm�i���o�(b�5t�&�V��$�M�C���#̢�!T ��9^�����a'��0/#LUN���Ε�n�U���c��p�}K�h,S��l���� ֏d`Oj1����T����

�&�����0�ܵB��o�b��o���B���wPSa�߳���kM mDk�e��N)�e���޺e��-��n획y��҈?rx�ĸ6�I��Z��ّ�]�Wځ�c\<f�7A��
��u�b���#��c$�Q
�Gw��,�	����oE�hB�"7�rjdb����e�~���_p��Go���'�Wڼ���{��*������pq�~/[��_�+��038I?�L⻔��W�0R�3Y^�ű0����@Q�yy�1A���1lք9����������^! 0�ϮQ6�ͺP���8�F���u[JF)�67�o+Ha�ȋ�U����	�l�Q���q?�����/�R�%PrI�#��otx!�3]�4~�qpW} z����83���k�7����q�=w����o(Ɨ��8�Ԯ�'��n��U�n���t_��X-7�GG�=�h��or�]dS��V{w-$0˰�Dx��q���/
�J�IR�AP������F��P�q=q�o�mu�|�7�|���NeIC��܊�.�iȉ*,#D�����2�C��#:\��3��m	^xH�4�^�D聉I��kI��B�Ձ�2#�OB-<�
���~/V��դ&&��PG�M4�δOֈح^&��.�\��U0���ת����ք껓\�=�K�j����/c�tu�B?�8�M�h=[WV�rvP8;&�`�k~K!.��%�b�Ss�&��E�Lg;�T�2�L�+R���ڇ�5���絛���@�ͩ]����ʀ>���"����c��Q�N��ʧEuK���PKF��rߠ?�xܰ�65"m
CQB�ȸ�k'��݊;���jë���N�)�H�%�鑹��t"~�X���T�(�%�堭�� c���	PKiu)���ߺ��J�:YX��敕xT�c� ��$\}�x�Ӗ�4�G�*v(P�v6<샭4O�r��+䅵���	��c�Z��z�D?5W��K��,���4��%Y���3�����E���}�z��[{#ɔw,�*�������؞"Όmv��Y؈����~�ah���$�&�A��_�b�6�Π�Jd=$G��፵Xb9%�hv�e�E�6�<a��>なP��ܐ��|~;��P4T�:>Z�6D ͉�a(�2�����Jv�p�B-���Jp�{�.3^�Pg��5��@z��#�ǢN�"�~��1��L��c��*$��?HS��o�?u%�C*a1q@9�O���B�1��>�p�|�(�ts���f)�k�!�*u�]S
R�9u5�0հ�Wh�Fr�=����Q0}����c
NזS��7�[0��xNؠ�oZL��)+�,9d$M��/�f7�	��xE��xe���/��Q)iR�#�Xdj=3U��ՕJ��\����_(����J����C�5x�Gg���N��U�`Q��ضQt9\s4X�*)��p�ߒ��n-y�>?X H4�_+e��GU�4��5��	��J�~�u�Ȼgv�B#F�F�1���R����jy=�>H(�!J��L�2��@z+XS�Jʻ�T�Rh���5By�����ͻD��L���� �i䑅���_OB���g�:�*�%( �����YiΔv
��6��k�����u��]�R�S�!�ӌ+S1�e�䰆�Q���V^�A��ȵ���K��ɖ�`��^�׀O�\��
P�����٬��&�/򫟆�-�s#/��$`1a��y�T��Ee_Ӎ� ��^�����࿇-͝,�c��;������Wn��|' �'?�,<)�,������`�9̲�����w��O�.S6-��[�C�������s�ټ����۔����{�_>�ւ�٢b�M�����hl��ۃ�xt�A�8O��[N�|�5*��`p�q��p����
���v�
�m<iv@��u����d����o+��IP��M�g�w^�#l`l/TP����n�#/W�i�:�Qu�`�oė���T�?�C�j��6@8����:6��my���uD�Q�����Ⱦ?�1��V�ԝ����ư���Q?W��OmP޹���oб��ej�̜��Q�>�U1�?b<��y����r�e�l�+��ͪ-�@��0�(���@6�~�Qg6����>Sѩ�VrUV�k��2�XJ3�o�;2W:�j�11�-*��Խt,Ff���~�y}�K�E��d3~�&[[[L�Cm�B�Ad�H���v,9 (�!��{a]�]����(�vs��z*�iCL�ĉ���(��9bM����qn>zi%����
�ϕXjxdG^$�Q�<.�U	=��.����i����KhAZz{�=
&�����p�(v�K� Qd�}G��~��}d�?�>�S�a{��^|}�>�#�ұV����m�e�1�6
	����3�\�Za/��)E�w�sr��+�O�\��z1���� �u	5�D�f-gm���Ե�k!ݸ��@�@��Z�4<iy�2׮M�p�W.�DL�AQ@߈i���3�LѦ���[#L����+@����;A�NmPK�Y�,�Ģ*H�XH[�<Ό��:'�P{"rݒ7�6$q�À� NK�`�v�ư�[�����WF����l�?�@�?�6�K�-#o4���Kn�<�h���W �m�]Ph���d;f��&/pe�+���!S8V6��[.���B(�����?ԅ8�+<e�`r�d[�����&MC�Gv���Q�X�&27�/#U�E=Ґz71ik#G�WmH���V��M����п��[���zgV�Ω#�]Z<��$�F��`��2^z��Ė�p�UHU	PlB��w�)E��߀9Kc'A����c�6�������$�Z��LHJ��l
�6u�r�[K���y���
1�W4����`m�:��]��-�����|�;��,L�G�*|-$�����i�r�6_����}����?�Of7R�\��.��)��t[��7�$nd����\�V�����XĂg	}u�NW�W���� �Yo?�
��:�腆k��v|���- �0��z���*���IQS�O�tg��'O:į0Ap��@������'�P����~TD�#Sŀ�k��� <�ۉ}�4�
.�nkjz��]�����~P;��RK`u��Ѽe�K�J���a�b�)C"�b��p������Y���M���[3������h��K�UXXJL4�)��媟�d�Ƿ�\	J�+���l������Xf%�t�&ܩW���U�k��6�|��%�Jo�JO�L V�:%�����@�L,���2�vNef��#����5j���vC�[��J��e���<�����V�*��ML�ϼ����+LSWn��%#z�����Zo�	�]�ލw��k�䁋"�ƕ�d0�7ޮZ����̂R�d��{Jq�ez�m�g�c�����=:>�Y�����)�Oz���n�	����i���x�F8<����Z;����?�'U�^�s�,�p�,KR�߶�C���)[w�:�V˿��9�>�Ӟ1�2Qз9nS��6fKǇ�5��Ł/�<,V*�)�cK�t�F�jO����Eq �6��#�1_BV(�\L=�*^O�\{H)��[���Beʋ���Ji@�~x�����R�7qA�#��5-��0�����#E�����R^����[��Ȼ�'Ppu:V�"	�;�^��[��	=@�*�G-����E�]�2x�:~t�\MP��ѫ�F=P�.�Q�j�q��܅DS�3��{b�⚏7A*���:��y3*v�U�Ӑ<�X���"�I��㾌Z��c�z��Nuzkw��%���"~�2��揉D1{/��&Ь����p9��i2*韓,J�pL�'�L��mM�.4�J�҅���/���jv���Ȯn��£h��4��,x�@:_��J������]ZGK����R��vzo5�y$�&�t�?K�LX����/�8��h�!�[i�hi[�}[PH�E6�m���.m��Kn�͖L�����K�����Śѕ���a����w�[mY��5�ɸpX�6���f>���ڇ�����?MXzy���%�J46���>i�]���,���ucU[J	߹ܪ3iD���% �:H]�;>�vN9G��ʽ��(�HnE����V,�����gY��f��1���1x]c.r�ҧ=UOr���[�)`�u�y�|�ЌL�ض��12]�ȗ���p����;�zN����
K��Z�� �l�%�֦D�^��|�r-@���I��z0JR�G�|?a>u�5�21J�L�.<�F�b����8D��c����͐:2#�ܩ+i_��t��A�?��ӻ��H��	w]t����eH�;\�)M���M�_`����i���9Vt7r,	�Lj��Z�C���v<#T�+~o7b�ܫ}��({�T�fY��$�pU��>���� дd;J'�O��:\E��䖯-	�5�*����KX:��9`����R��k��|Q�#��_w&��<3��ɽ+V��G��&
S�B]+{Hr	*S^�l���Eƃ̱Z/ctO�К���'g�,�8�`-E�r�Z �aA}h&H%�,�ąy6�P�g��e��/צ�O��� ����#7��Z »����GZ�"�Oy[v��:˪_Pz��t��kR3�_#�{��i��x�h�&�N�po��9T���q��P���,�u��cs(�Z	8�%��gZ�i��}55�'}Rf�5�)�b�RV�ӡjs�@�~���Zx�x�WZ��̙HL4��87�13]�q��lK:�ͶN(��J�u��#5g��6:��>��]�Э�Sa]�;��E�:�bg���рт˾a���v�[���^ -��:��p�H�� �|���(�c�C>�15pf��X�ai��㇜�J	�v[������Yf�b�l"|;�:�s�
5�r��,�����dP��g�������w�R��xR�I=ґטS�=VAg����"/y�1�M��N�Ie��� ��j�ft�K#Q<n8�,ώD6��%�~��xL���K��d��~�I��:�y}�H�-��!��w<=x�@\(ZY�7	�h�XG�˧�y<Q���^�(�OX^���E�$�E|x);c�1Xa�"_r��1[h�y�¿�
_�%��E�f۬9��+I  {�wk�7y1��q�e�E�>^r�
�P���(�F6�q�x��(�55J��m�_��������/����h��� ���f��%T��ݐv�r�e�[Wr��[�t��=�r��
8�'
R�Y��\@?�:bG�S���_��Y�p��.�h����&�},�b(f�ζ��W���D�'낍gT,��?G��C<ygٚ�;�����Li����G2I�7�lT?���/� �D��#���x[��rt���G���n��&tY{f��w��o\g?� < �I�Jcw�B>x6�Lε���_�FS������<�o��T��T�3\H�����l��&�_b�k��N	�OGEb�L�-�M�P�vV��-*+������8��ޘ�ߊ��@�s�ُ�
����Ŭ#8��<>��vv��W�K�;��a� 0��ZϏ0����¥x���/��z�|�(�o�(J"�w=�`z�2X/C�[�Ծ�DL=���U�-�F[��UG��b���(̟�����@�M��~�c��iHA^MI�cX�vn�4�*v�ٹ�1�.L��)i���4�n�mPv���ftg�@��jsW񨤴�\��P2��#�Mc2��j����g�k��0�Ġ�pe�R��E�*�2�In*]���q�QA�HOI#��>���n���bNV~7�,��Y�g�{U����Og�mz�&}JK���Z�������/�g�N�-ܻƆI!ZT����Z��i`�Y7D`MTqF�U�{��5��
l]HUޮ�B�^6��ܯ�o��L��LzP5�]� ��ho��QސY����_C����;�Z]7 4�nҔe$tw�g�)�������������!����m�*D�Se�a1W�p0�h�_��� a�r#Z��=��}�����zB���M��-:���M��Ufu�Hع��z(����f���4zu��o0�ڴ<o��.�����N2)��ɀ��r�
;���P4\���[��X�v��T��;�j���<�����T8��̽���|[U�5�R8D5x2�LR�ׅ�.���J@3��P�Jf��qmI��YQ���p
$g��Dp�jj���gu@���γ�*�(a�_~�cM�!�6���5���ӷ*B� �t�ib.aɮ��	|z6�j���C�~�jͭ���3�gF�l$ ��p@���H/��~��X��tN��zb�_}���@ɲ��4��bJ�*�۽QЌc6ؓ>jE�7���;g��d�d�^Y�O!H�?$P�~�O4as7������5�v7�nq�O�����#�tt������=f�X�&_�9_���[�6,�>������Eb U�U+rˈ
�UG+SXK�i���h<=�	��r�=>���]>��+��n:~_�H^��Q���sn�+,ۻ�PTʂRZ���u�7������#�����&��.t`���ơ7��Ϥ�V&��r�jf�&g�;�/k�C�r5�Ǌ���[�+�μ=���N@�b��#�e���+:���unz�!��VWbgW�#�4���N�o��l
�%p��z0���-B�=�խ����q��^���rO����[��0�[:�u��Ӛ�-a֘G8�%f�ÁE��M����~!Co�1�=��sfa!7����Z.���^�J|��hfh=�0x������,�mU܀{osRV���N;���g�	8����_�;%`2'[��P��%�2�� ӽ��/���WOJ��)��#��o��5^0j%e�� j,J|I��9��[�>�>� 
�G�Qy=b����b�#)	��H1En���Q|y���60��>��:F����u��d�n��x�z��z��#�{?m�?�F��H�$��z�6����l�x\��GS6��*�:���EgC�e�Лc�'y�j��P�n�}� m1�G4u�v�4�,�X�Px��]�7�<1�ߛI��m��)�2�����$��p;.�0��5�Dݰ+<�A~UYx%������g"K�ݼ�_���"p�?N=�x����N!�;��o����?��9q64(�%B2�23D�����#BPC����,b�~���b2"�v��W��ǆ6�*��A�!�٩����l<��V�,� L��¡̀��@%���=Z���<��}?����+7�0_����R�M$�婀/�$�W��FqeA��Y��l�I�T1��5~�엥�����>�J�c@S8�y���f~qQ>x���8��lՙ�@Ĥ��-�O��A'�c�2��-�/��	�"83S
\>ﳷ R�mv�\�'G��HI��������@y��؆�w.A!lK6���&+��i��4�([a�"l	tj�!���(���2{K
�P`S��IP����O��!��b`�pI?�r�X���,����6�'�bIZ�����r`V>D>{!v��Bgq�B� �ԝ6e�'��_TE&�>�$tS���MN�o�$4W:���<<hK0����,VQ���7�_�Z��[4l������Ҏ���o�v�;��{��K�y�r* i���dA���C ���UF�7a
�+��*
�'����n5�ѶUK�h ��_�uz�}�N	W�7t?Yf����F?�>��w�UE�۵b�H��Ԡ��];?����8X_����(����2 ��/�n|��U��K����=J|�;2(��a wk���F�i�rR��b�:C���8�Ӂwa�Fr_���3��N�(i�q�f�W���G��	6!�����rw�E/��l�]|��8���7`I��O�Q�#V)'�\?5H���Ң_.����Ĝ'W�Uw�<��r�m ����/*�)�08��{�U��(������ި��xlU`�3z^�B�bv��U�1;C!'yt����O2���z��-�?�(�ʙr�J�jw�]*� c�1����]�?e��](,Z�txrץ]b�dN��x8͢=�"Ǌ+G(#뎈�a��cR1��?�t��8D���{�1:�ͷ"/����F��A���Yno~!�6B�iFds"p����t��=%�uy�)CG�V����+��j���*y�B�a�w����zNr��
^]wMiWp�������ch*�z���16�bS��iZ]DYWZ朹�"�q0�mCr�s�U����z��xpl*��2�;S믷z����h�p:ٴ��;_v��j'�?R���,Y)m:�uJ���_��#��r9��cMR�
�B�(7O#�xG�T������>
�d��zvU,�G�xQڱ4
%*���Y���$w۬h���CF_������-	���u5/�J���y#����7P�a�H�!��g�u��L?A2�n�h(x�٭�
a����k����&�dQ�&���.���Q��eg� ���x���M>���G�"/xƢ�#�_vmS4�X��ݞ�ꗄ�Α�ɛp>Ƞ���D�������`�\�q&�1qA��)t��%9��K�j�X�{rIWf�py]Wt۴͔�O>��ʅ�/t����f�;&���C��JKJ��l�]>�r���k
|����\���_�U@q�<���>�մ�dZǗQފ:z=0�,4P������x,��nj�}5)�ㄗ�e�� ��8pꌻ���	$[$��:���O���l���X��O�=ER��cч�[8a(Sk� ��8��=~[�5��ˇd8Yc*������VH��9��h;��_��r��L��tڤՠ3vc?c�5{��-�ꔫ�
��篙�!q/n����,�����F��%�
��jG�$��,ax�Y
����f�M��m��;�b�}f�5�c8�2(�/���߶������
w�`6�����2:f�[�قb���Ia�b>�v3��F{x��D��Ա�ku���"�՚�H��*�G�e�o�d^W8���Lw���AP�u���@ m��$�� $q�h�vh�f���a}�	���]#*�w��w%Z�m�0�ŎN�{�]�}�m}��^�'�T�����(���0!N�bn���TE�f/����#�P���ԏ^PQ.�-Z\���F$�%n�Z�׽^nlxlB�Gu>�v5�1OIptq=� j@�~Se���Q�^t����?�����-�d'DE�;�S�fUK^�;�i�B� ��Q���`�G�N�K7^z��A�A{�8���U�2�J��٫K=\��I�Y��mP���N6\����*�<mɹ�A�Z�%0���:Z�B�H-C\�˨ �eК���<�:J�N�s(��Eأ�ȀGL���k�w��t_g"�N.�f#D�V]@��6���!O���+lk�A��� �%Bk0�l�H�d5A�W��y��{�ǼL�A�����/����b��
��� 5�r�ej|�m�<����dh���[���ä�Qh�!ݍÁE12;�W�ޫupƓ�$���[K�eːa�*d���[^D�0�����}`�{H)96���R��oX�1��ܢ����t���S�A�/>q�X\�0�"]T�l U�Z�!�Š�+�R�#"��[��Q>m 5�d֍S����ޒ��@�4�%���AA)��oT(9j����vh�[���B�7Q��0!�rR���(��>���@E��b�X.�C�u�(Dԑz�Q�"ӵ�97�[Ka�ioyrb���]��*���)@ꚰ����P9�`P�L8�P�]�ٸ�����B6x�n�o'�K�ҷ���4�T��P�������s�E� ��pf�f�~٥Ksr[�@�^�
�ʱ�	&��Z]C8�t~Dw2�,�{&V�1��#�_ۇ0�Q�9-�� o��mr14�+&�jn�%���h���7��%���43�B�����z�N7hf�~r���2{n�n{Ӏ#�;����5���B0o� i�./��-�u~>Be_E0���M�b�)¯�mf$�o��aDT�.�Ya���Y����#S-e0PD���X7Ɋ�5��L��&�-����^8=�zI%[Lc��}W�{�;~W�0+JGV�Ԓ�d�o�KP��~f~Wđ����LB���C�}8��L���),�dl�b�ׯL�6Gh�g����Q߻��욻��쐖7��Y�-���ё��Sq6c��Aؘ@�m��0=RN4k�?~nZ�%@��t�-�K+�z""?)�b��	Y!��2��0eɉ�iՌ���γ���2�Rn�Z�Cg�s��)��ޒ\���p��<�p�#�X�е9%+�ʊ��"�ut�9���V�N*��r�T!)SB��d�L��p]w��"Ȧ��p`器E�������0�\ˠ�	J�}K����|(��)4���F�H�Ծ8���?C�rT�U��3Y�"A���t!ᚶ�[���^o��P��8Fom�������� ?�U�Hu;7S��M^)�6W��p�" ����P��VH��G�,t��Tm�p�����$��i�(W�N��7��x�R;�o����ى�\]��ƍ�������B��M� W��y�=�ٜzr=�"Y@(�mI ��C�@��$��=���ʀ�ٙ<^��K��Aٍ	���N�m4uvpbq�7����J���@�Ut&J��u�ݤ[�/Tݪ���f����P	��r,���i�t�\Ԍ�Mʑ��c<k{��tOX��(9��I��?-U���Ճr9q���I�<x��
 ��(�Ԛ<�itj>�?�>��x$��=�@�
�)�>"MT�f����]BjC��i���}�^�j`qB�r�����y�sX�J贈�X'%�DҶP�P���s]H�fI��I�r��- )e�F1c�<�t��x��H�.r�z����31�����Ͽ��Km��p6E����@���1F�C끖�=��n2�ԳC�ڠ��[3h�d�y|^���]$��(��H���bC�n̂��h���f0� �k̖�*DZk��}�)O������Qv���L6G�h�DI�x�V���2���������z�*#OI
f�i`A�놹�F�9�y<�!���}�T�"�HA���suX(Y�Ps"��V�_�+�F����K����F��{	��cg6�.�S��j��Z�@Nާ�� ��;��`��[5N��|�����if���Tͼ�"N��x�	�����2\+�`,W��FxK0U�X�̻�>ԓ����)c�a��O�v#\!�����'��4���k�j�Tə�˙�NI�6?n�.{kH�Zœ���1�	���~�#{e�gra��L���v^(��[E++a�8�g�!e���qryi�ܨ����ι���DZ��\�*�E$�z�*���|.�Y��IK�ـ��Tωz��lYp�Gm"#A7t�b,#�������NVd䩵�jz�&���]7��7P�Ӕ_'�3�܀΄����xR5�"d�
�yKRc܅
����;g�Ѿ����!|N�ʑ��
A��4؉f=�!�ӖyW:_sn���1��eRx�F���f��-�ۛFg;՚�
�J��n���k�v��1��HƟ��?�<g�ϱ"�*�X��3ͱHbpt[WR�%=|њ8�x�+��n���*�G�C��ؓ��N+�e ��d�##4�A�&uP7�rj�t��21ܘ��'�`|�o�HJ�Q��y�F��y�T�����c�Qn��C>l��9#��g�j�b�������j��&�ZUI��e�O)Bc�%��]2P*���a�#�F5��%t`��	�8dee���WKw�*���>i�>Vz2������ơ濊<6�L
���Ch�?�8���;sD�\�8ɮ���"~� ��zg/'��0-`G������'��r�g2�#%�!��.�1^nJ���\F�xD*	�W���AWq�bMޜ�^��U8gef�qmo�m�?.���Ca��vE�7���8N!�O���OM��i玻/|e-pQ�.��^ ;r!�yW�I2���.u$�F	\�k�q���Gi!m����20����`������'��<y'�bF�/��47`��\�+��1�/�,Z!~��叒��U���])@T<��L��/|�c
�[�Cake����m��(qõ
����|I{���|��u;�O�(��}"�������YJk�NL��Dx�\�mFliHN�w��� �S�#Р��{�.
R������xn��D�0oP���@���N-�ȼ�/�+Q���L����1mSr�%���
���r4¢�b�Vri���Y1tY�M�������4�{*�]h�6�A�եS.���f�� Y隸�kC�Lj��p���I��Q��}t3zLW�zw@���L���ZW1��O���ď+����.���x���A泖�߯���_U���ő���B
ْP�*vZ*�8ھh8�RCOH�w��쮱F��E7(0+���@��2�FO\�`nh(�э��
�� �/�)��QP�����E�@{����'Z�l���j.�.��y7��Q�3AE���4{d״�|������RŲ�ܱVʽvr�mMÜi,�y�)j���M��b�	r�<��$��1��CX��D6J�PF��s��A];ߏ�aU=�ϒ�����0�i!�}:�W4�:�ZI�<|'.1HX(v�i��� m�W*�v��qnW���M0�)�Ȇ������'`a����V��S�l���M��ܞ�t8���)����T�I�tb���^�B���3O*� �d��c 7g��7����3���0�WN�n��O��4| fvD�&�ܵ=1��ky���1�	w�qx]�D��Ԃ+�U�t&8���;���}Qx��h�Y�_���
@h\�6��8�;A�?U�0������u��E�Q�`\��X���Q����V (�&3�ji�U�ѿ1W�|�{�)��'��D7�+'�����qr��W�}����1�r΀OT�T;<2NٓN7\4��k�<��m���Xݡ]�S��Bu�n��C�g��8�Va1�(������>&��? ��Oi0S
ֆ��Ͱ�+����[=X��k�h9 9�UL�u��b�����l�����B�a��;ε����Kh	�`�ꉳ��C#��q��.V����icс~IG3y�l� ٿ���e�H�
��<Vp�ū���yv�D�%�t���o���i�-,����ub�v�������:E��K������a�yO�C���K6=I�ޓ�{�y���)�7V[�=�Z��[�=_�έ��n��)�|CB��?<!�&�����WKQR��T�
9��W�rWQD�fPX�W)�Y�V��s������
H#�ß���E�,���ј�z�P�zg
��!>�B�\�N||at�D�E��9[OOW^@iH��,4#��tHb���]$w�X\)��e,6��]Rrʶ��!gΓOw��7~q7a�8�,Jwk.QϔyD3O��_�A ��9
�)��?'�ʨWc�b��Q��t������5�n��O�¤X��1F�I_/ʏ�0Ӊ�޵r{�=�ωv��咰��N_�nW<�+˥[	��A]Y�W稻}��2������ �x"�8!4����*v�8}��?SOM��I��b"C9��A_��%���8.�-�7I�l�Ŏ�����`�����E�)b-P��@���� ᥘx�������a��oı�9e�ܒ���5xo!94���ӄ�e�NxJlP:���K(1����W(��(<�N��{��~�n,��Vsn�ch'k�SY5�Fd�1� _m��A;��LN�u�
���\4�<�/a$3�D���2b��[x���; i-�ek?Ӄ�-�6_ �e!� %��4!f��zzW9�6arɒf�?�!27�E�5��
��b� q2�([N�c����	�����*���_6@���-V�[�'�x�``��_���W��#��Zҟ����5U&���	���-H�CwF&r��BߢWu�T��r�Z��	�Rq���69Ka`���*+'W�a��M����u��n*I��+A��~���3!/�!�� ʋ�ٓ�	�w:S�$�P6��
T������8h�Sc'S��Ө���1h�{��b8��A�!u'�o��Qc,�癰��n�#���f�5`Ta�Jƃ���RӱŃZ�Tg�]V-pȝ�1v.~�h�@%�zw�G� Me�툢�r��G��7ؤ\��N�l���h<�s*n%�P=Ĥ�7T8;9D�m�1~]�bD��F�#��q_�G�M��?d��>:XD$��-��q�m��nTqñ�/mB�l�܆�G_=�H���wy���qoD���7T�'�|Q5��g��%"�����&��q��`��66�9�ψͬ
H!����B��)m��z�����ޭ���O��o(Q:�%zd�����i�d�N����"���79,v/a'8�?��;�d;k=�Z��ՀhB���j�n3��v�p�4��$��B`J�`םY�+�������N��a"�E2?%=>,�����ԂX�ɞ�����Uh�����d��o�#��ډr�Oz�x����i�S����`LJim���s��b���Zg��<�Fy�s"�P�l�ˏ�"��~�l����R��9|y�Z�;�N���շ������D_�>�}a��֗"�Vfά+�un�,���9����k���?��=v�%M���Q>��_��J�44GҎ^�0�O�TeFh����V=�R����'T�T�{0k�/]����0�I�)�#D���ͣ��儜Q_�12�$0^�ǅ�<�]�,�3VY$C���NrթV�Zhx@�<��3�2E<��4��'�C�W��,��E��w���o��q��L��<_�r�����dH�ȂXU����Y�k9�����Rx���Г?�����m]��Nvn��**G����W�9���M#[�&q�sD{��.&-��c��g��&��w����B��5�cA}�������E*}AO������+\�"4"��[j%�ce�A�jp�P���i���/�z�Y��N��'խIz_�8�����t�*�>��`�f@ ����
D�骁��+L	U����#�ͥ�,�V��n �:)�k�O�r��P�����P�4���Ͼ*Ȋh�c�ş�ac2�7��[���\C�O�@��cب�$zr�����J��&��,B�6m&�*4����FBU�����gi��3��[o���<�CM󔯐�W*���M��%�)��pF^%��������KAE��t�%�DS�����D�&�FQ4�J��z�{vu6M��ڟԖUS�h��Cc'z�A=���ۗs4��c2�.~\X�(G�*�h�����G��	���U�RY�����ȼ�#n/��LHA3��4�P3
�(��	� ��72��`��JL&~�����po���s�������l��>_��6�$�@ �x��Bp�v�9�SC
5�9K����#tG�_:�Q����f�X�E�aܖWc�6D��= ${!�M��ƌ V����KV�e������U����N�.�C+p�,x�Ox�~��9�����N�`�������(��L<��q���[[QV������<_��䙵x7�X�!PG�S�e?I ɵ�^j3{�|��	�
���+HK3j�׋��:m�M��	��A;ڸ
���5Q�@\a	{�|f���V��)���yS �Ҏ����D�o�`n����!rW��|ﾝ~ܵ�o�$�4�pT����6��	�S�Nfj�f��e7�]er��	�Tǯܾ:ՆN�rsV�u������t�湊Z,������SxYݻǀ0���B=j��i��>{��ڲ"�e:$���(m�n�W$�[��F�D�TJ_�m]��)^�͠�Q��u�a����Z?�Q�h"����2(*��k�3��"B�q�hʏ	^�eDjQQw���41��k���N;`��<��.,#a;K2�zܴ�V���luF(/�:��7�`� [;�Syj] }Xc�!��y��s�ߩ��C�u�@ �>4]d8 ��N=p��4��%i[rk������a&0F�4�x���qX$��B
3��,ޑ�񱒚t��[(`r���߄��B=���1�5?a��li��;+m����R�k{�Z�{<v�����4΍�gT�H��d9�L���=�������/z[�;�U�Z:Kt�	u<M���O4�~׍�E��$u��؏�n�`E�ᐍh"��
����"�<���ʜ�]X/q��V�a�Ǎ�)���=��I��P�[)��h^Abb"d����&^CD� '���9g��oN�Y�tsĈk�>RR^
�;��p���bN�1 p�Ha�E�V����f�u�Va�$!�lj8=����,՛�i�_w���C�q��V���]�#�[�ѬY�ںs`��)̍ƳhN�;t���W7_z_`��Nͻ&!�cznovC��%�U�,H��;�#�)Y�6栅�kj�\,l��z0Ʀ�(Q�p{2�29�K�CO�xց����~�a�O�JY��ilC�c�P%�M��ݽo1v����T�9!8�q�l���k��bw��l��Y�4����}�1{tTp������`nMjx{�����l.^�����hɋ�`d�)��HliM ��OS���i/��M��s���#����,�v�["��?4���w�� ���Wz��)����_��Ua4e5B��|g�!�] G�H���xbg��`lM�g0�X��Z�y�Q����ѹ��Ō
���r��3�"�~��x�A��ɯ�C�M,���I �~�������r�)��3c#|B_S�b/��dB���/�������V��%.�/@�Y���{���TFNx��'������rR�EڅX1�����(����ɣ6O[<�������b ���d���T���
�m�������YjiY��������ʆ��e����.��+ ���.�XVY�����7m��J�`5�M�y��<���a)Zjо���ٽ��Mձ�Qd{���9�%�m��?r��/�� *��89�?B���֛ٙ���1����WQ�J����4x���m2�e�	�	*_<F*���1D+ꨒ�-�G����]�&{���
�=�.K����Jzt)�PPT/2�R��q_#�f��0�)��nĄ��\9�$���j/]6��� k#�PĬ��W%�����<��{C�����H.ͥ]���Xٛjx_��?i��c^��b�#���c��r킗M���o�#��02�*Ty�z<�i�i��P_�l^���w��=�U�b�!yҟ�>&;�5?'�2}��w��+�����)�D��/p�~�1YE�"?�#r�kLpGK�s��:�7u/�!��qc;��L��h�D�>z1XV��0Q#8HtE�\ŁO�Gﯝ��<�?�)*���49 0q� ����ށ�Ť$�\���?��U~�m*�h�@���#����hW
p�K>���E�i�Ο��|	F���d�z�y�mzE������!��9T�щ�>fpBࢿ��>T��l�n�ASZ�Y/b�@��K��s�[XjJ��xAZ�W�)Ģ���o_��S@H4�x_��6jV��U⪂�vv�Վbr:�W@� d�	�&����bw)F�Lܵ�w��LSm�;3��2�}n�ֻ_�tTK�(���H�q���
�+�g���Mi���V.�i,�p�΁T�]3J�s�ϡ�dϪ&��K��ɸ�L�(���p�`%u����n���=�ga���q�kM8ƪ�,{9�ҁ<�X$�\w.$�i�Pь��;�W2ꀉ�"�x,mK�5�>N,���.i+9�k��p�7�����7�Mf�{����i|sYM͹Y���!y�4�߲)F�4p/��u�"��?�6�����t�_&�º�	��}٩vϡ�����Qӌ��ٝ��6럽F\��«A�i�V.��zC�����;Ƨ��5�$���\��Tp�����Ù�u���_��{�1/�%w�(v��yሩ�]�Cԯ�G�B�G?��ެ"�"��Vx�p��j�@����;��u��L̋A�D$M3n�"z	�&��e�v��`!�0D�d��J�çK��u�������`��y�I�vKn��Ǥ1L̅��r�TH�8^��`ΦK���w����x��x4��b�$x�>��o��Iљ��I�`"��kCy�� �F�C��u��$V�*�d�ʟ��i����4��6��T�]lO�9�+���,���C_������IY��'�Шevf���}�řJ��$�癞Q��-}�Y�#�:��Loo��r�8�H�X/�23�=Ԉ�"�����p�qۄ��A���![icDh�?o�6���͖�4�];��T�#�6�N��A@��m�Fp��EP9����ln����5f�Rܛ��%Tb��5��k��p��R�0�p��x�8"6�V>Fl#̠�k���.���� p[teG�����S�\�"��0O7�7��`�{��Ŀ���?�	I�����6���0(���*p��4#�z�:TD���l�)y�<�I�_rWfӊ9&�o.Hp��4���et���+��(n�j;��g��$�w��y����.i�v*��1u<�V4�������W�'��������/��3����h��7!z���E�~���0T}]�yA�P-�c��*�$�P�U�����5�3w����%�d����o� ���	��R���g6HķVs���y���3�j�ek�8���S��	o���r*��E����?v��X�4�k�OIKi�x�Ȩ�H�M(f�߫/��\i�h��#v�Ú���/ڏ̛ȶ�ݹ��9�q�N�{�#%-�о'�]�2��vu��7���0+N�4�E����8r�ԬP�
b�5�1[����4�qO1 �m�
�;$�'�h��a��<���k����(��LD�م�dw�_�zݿ���@&p���
�_������9�f�Ǻ�y�?B���4���1[�sG­b�$ �����:@^�s��Eb
4x�sDс�ٺ�V����E�,�;�%A��,QX����(Lq��>Bz}c��ݲ8�� oPLf�7dF��Vs8āL�\��+O`�>dU.��z��Q��.#7K68	�
�ѓS`�~ ��RQj|�7��7	a0�����m����L@�f���]�|p|������ J8��c��x�]�/0�t	�.0����1�_�0 �a��F��p-p���n�^�+8Ei�U.1qo�$�m��1XCs��� r���]C�$�]�I&HE��i��^D��N�����(��!������H|���]�ŀ��t��xqw'�����53�n�+C��R���tY沗���ߍ�����pS$uQE.��we��x��jR����{��*+7� �C�
8Z�����R�=��9Ro�]�CסZڴi�Wv��>Z���*�����5���J*��	���l�����v6�<�x��\W�D���|+�7:>Gr�@o�f��6K�NG��o�K�zZr
��!�����i7Dƞ{�����;����ky��G�]�S���I�Ӗ�-�*^W#�q���G�Ɉ��|��cl�$�l�PX��I�puGI�%|n�e�dCh�
�j;�!��$�I6Z��"Q�*�C�w]�v��|�����C�=�7|M�d�7I-��'����N~�`�;���J��=�o:��b3�����2O荅ޖ��\|·�l��_�j��c	h,�C6d�9QS4�/�WH�����/�s`�����=0�A�eX8v9�ݝ�e���(O���o�MX�Vn�z��]1UNN�9<���Bd����j-��l/�^�#��zx���gXgy��	�/#�(�Ɍ<��u�]�(�٥�p�Q�?�{�8���%#���8���5X�>�i�o���V�O���O��L�AM ���ߖt/�,��X[23a�"�Ԩ�(Mf���ӳ����:�����m[W�]i���� ���/����)��[���I��Tx;#�� -�Q�����S^�#���YU?F�&�Nd�eH���!fa#���k��#C	��ؒ�VT�u�r����ה����3 �u�2��w�����lTt���̊r��LI�{KÑ��LI ����`�d�R�V���B>�ji��t���+�5�C�_t���ľV�PB��Pg���oz�h��O����G�9&�.>O��m��y·*����l#|�;}VJu��uK[��>�h���W2F��.Ihˆ�cI� 
H�9�G�������X�@/z���]���w'���Ɲ̆ۛ����{��������������P�������G�r�UIS$�_�t�U�@��s7��u�%���#f�*��3q�o�\��`I^��Yj�X�E/AcN��,�̓��j3}^����y���Adp���r\y,':�޾U�얳v�S�?�%��L&��s�W��E�Q�3J/�m0	��1���AwY32�BX3�I(� �1�\8
qЪٱ�6�d@�%P�@���_-~E����r��oĈ���ګPNG��iuN�Y�ſ�O��Öw���_�t��._�����Q7O5D|||+���=�  �o�K������*�7*m%�'٩M����|�q��I}� �rճ�o�����"��D��T	3�r�}�@C�%���n��9d (a�?B���5�HU�嬽��9�S�5ۦ� ;�ӧD]�!s��c�rS3m���O���"���RA�֋kh���	Ϸ�>װ�'z�p��'j~�1Crm38�˓��U��*!9C;�����������A�i��w���i��_@��T�j���Q���&"-J���C���N�M����X���X0C�c�q�-1�	�騠�S�5�.`[|�ZV'	>O���D���V.��9��^^�֜�� )�f��I��YK�p�
� l(-\�W�%�%[A9l����!�qAQ�vvS���z���C9s�5]՗r�Cr2+�.m�����q�]'�S��u����wg��H�jO%���Pߴ��P���JN�����d�����A��7�.��x�[���o�E��A>!�\s�C��Z�Z꼩��@~��vj�.=����k79�N����D!>iN1��� @Щ�>8���]}����B�$b��(�����$�mbZ(��o�-Ko���U�H}���Ohq�ETw�ePk�/�����ީ�>�1[�ƶ�N�l�b��N��z(hB��8����J�v���ѧ�5�����pi֒#���`�΢�.	]P�����T[0}/*�q��&��0�r��U�A�k�0Z6���d��|i�i�H��'N�2}6��G�c.��u�a��},�Ui/)L��:7��#�A�||��40)jӺ�p�ǇC��0M��9�"2��HBx��ozP1�c՜�qn��� �_�����]+h�Fxl<y��RT^���"��ty2cܼ?��3nx���30.��O�%_������d���!�ejomD�}Vv�Sf����V}0|ޤ���n;d�s���u��71s��th��W� ��5	~QPa���S%�/5[��[�����,;,Zy�I��}����$P њ�Ħ�������O��VنGP$���+3�0����� ,h��I��w� [a�Z�*;f�1�K�����qg��\Q9�,�bk*Y�
|�;��J�������r��ū�.��K��\aB�,4�T8���pL��:���h!�K����ܮ�I�(��Ik�j�y��Kz ��^��sܕ��E�,�9n�����q�3l%#�*�QQ֞tj���O��Ԗx?�sd>ӑPՏ�x���W���Ed
b�a�'MQ�{0N�N�Ȑ���\!�٢��2I�ׂc�D����ŶdQ�f��=T�+k�)�z/��0E�%v9i�ޠ�Z�*ĭ����Q���-�a-�'n���6#�R�!����qh�0��˹� K �w�1?L"�K�f.6_�eH�T���h�D�XU�U��Ff�$Y��.Muo5�Zؿ�]RP�'�N����S���-b����V�G��6m�A��b��	s��r8g.���ػ���B���)�w��J����/j�Y�d%-�R��<�����T��sN��A�<�j:�b��T��T�Z��	k&�,5�}���r���]\49��l��&Mo���O�����O�DV���-�5@���޾L����bs�ّJ����H*kgL��1�3�L>��!�wm�� 	�0@*q�������1�F�ګ���u�>��-�d���Ɩ	���0x�!3�(����1M{)c#Sa��v-)bq[$R�����rs�3�߁��j\L&�@�P��#��S�
d��L5���O����K���C�7wK�I�M_��M7���R�`�_7
���
X@��[Ζ�LR�����8�6����X)�&����@�Р�n�IQ+ ъ^�����L[ݩ�>yU0���F95C#����˄�.�)��EN�nc׋C�(l�4��jA��~[q	��9�_���t#]���L���R���GJ\�Ŵ�Ѥin��
�\[��ѧ�$�8� t��exӶ�`���
u��2!�_q�=@��P�c��׉�rŤ��&�Sz�/em�_��/7��ʟ��ى1��b!7"훆�8Q%��v�S����A:ĩ޸k]�#>ڞ��Im���_�N7��uX}SRG3�
�p�x�"� ����	)���Q��s�WɌ��$�.�A1�<�X	~��RӠ����8S�ڝ�����y��q�w��S� 1&�5�	P�ld^�n:���+Ȫ�@4'J�?\1p�'��"�Ch�3�������KJ <�F0D���_|�ޝ;8s��X����1��qW��Gd���<n�PJ�2�R���D��Xv����0�݂��.���\��]O5e3@�cl��^���N�;�*	1��^|�:x�^����MU����� p)���I�,�_���XQ��E��b��������4\��	��L�.�����r�%7�!eKl+q�p���1tP	�s�ln��g��X�z�.�sPS3� ��1����o�yt�!����2�~e�pTS��(�)���x깬����U�%t�;�x\f�)���K!Hg�� ��c��>����3z-N^�=i�KîBჲԭj.��6L��fJp�$%D��r�����{ZA��.�����a>�F�7ګ�|]��.�E���O���48о�30�� y&�>�����/KN�j$�P8���$���-_�H�9֡�هa=!��h1y��K|=0�~+g��$X�y�+��@)���C)���Y�OXmD��&:<�e�V�m|�������b�M(!�{�F%㲺�����nRݸ?	
�˛7*����j4�-��ϊi/���`����t�, |Hjs(��f"h�����G�����������xW����Si}&�,q�f_Qf�<���8?(a�G���n��ĭ��:%iӫ���T!����N�������|u�;TU����� pR�١�2O!
~��+����W�	�	���>?�|�/]�_Ʋ�ab��A�I���)o8y��((�Ǩ_^BҲ�ĳ�Ž�PyF� �e�U�g���$}��Zf�S?�=�h�� 3�9��5�Po�f�Z{Q=Zp�l"��0P
J��C�̎�p ^�p/�����̌�\9v��U�����+�#�o5��
��S`'r��ԫ�u��1Z�S���r;��-�d1�rA�égV�O���h�D��	��Y��q��H�E�<�n5T��+��LaW����[�Hv����=�*~�Q��ކ^�יv�\
9poŕՄί'鬥х�a�V)�먼�D2�z[t�.���g�d��ZWW���k��X������q��$赙�z/�� W�� ����rW���!���<��40�
_ǜV-YU�۞�1�C�D��8>J�r��"�.2 hm�s�x�җ��,qsf�,�G�R�B@h�R�+'5��`�r��qڳ[F��x��=牦�Z��S�� 3umX�s��V�#x=je���a���T�o�%4[.D�+X� �C�Tߗ��l�"��i����?��oVO����tO��w�m9<��$Ccg���7@@%6���׆�:�I�Z[�}у"��a��bEb�U��@_n���rra9�۱µz���/GT
X���vD0-�s}=�J��>���m�W�I�pn�^�.w���H����H?�*���,jA�aﯺd����W=�嵉�[������	\#X�q�&�`	2��W=��`���%8��oo�_c �<�&�В���	���@R�1!j�����֏]���>�x���clUr�G%.4�����ލ?��|>�Y�<�JL���U�r�\@N�} kB@�$Ua��:�:�S��$x5(���>l�r{���kdÄ�o��&H��4��Wr�]����s�U�jx[��2d}v!���N|=����r1�5Ag��=�����b(-�4J]$�}��[N���h5��0{�	���g���6��J��>�a�L�h$E�ML���}g��7q��ŋu��+K�fe��� ^�����8�CXL/ q�{x�,i���$p��2-��r#G�d)�~bn����M���(��tC���	�<_m]��(�>U9F���ohgR'��0�}��(��-j
��i�E��u��]��=U� zų�{�B�En�%���g(���9��2���2��9����W)2�� I�ˍ
3I�|�n�H��vp�ޗ��.UX�����j��^���y-2���<����sY-��B�E�f��?_O���L?�r��֥�u�����A�v�qg�������G�+\���X)s�	$��<R�f��\b�0b�A�A0�-�����6�Dd2��S���)X-l��	:^F�ĳ�����r���R�9~��~�ӂ˪�m���/e�1O:K���d�	�`�۳2d�G0%d��v�'�t]�1Kձ���_�����$l�A�k>�*��y���Fn.��௃l�`�.#Z��V��5��gZ��}���)uԲѺ5BB�$�U�g3�����pt����{-_\5!Y��5�*�T��A?n>����L:O�[�Vd�P/^M(rI���J^:���N��$3*��T���~���C%����"g3X��{�O@��C���]�LHCG�~�	:���('J̫X
N�G���k)w�i��� �2��i	����8OB�g��;���jp����{d:D*6����>3�dtV[bs���n�� �ID�|G�.��ID[·ʶ��j1�.�Ĺ�|��yB���Eg@� *���-�f�;�zZ��Q��l���闢�X�$�R'F�{�����'9��mo���'՘�*��Ae��P�.���gTs��1�&���9[�	��<*g!�i��+�g�E���{�Vn�ɺ���5|Do$)x5��A<Z#P)<�ĭ�o��:�Rzպ25@��°� ���C���+I��mjH3�X�,o�&
8�c/���
���]�v�\���)OϿ��:�� ���'��.<��F���r���\(��H]��M��K�	�!ߞ��k|X�V�m����4Y��SZCnX[�!�݈G�7�]\^��>����[��8m���1�̬��k��_J�Y kB�{j�@���ٷ�������H�nj7OF��[ْ�s�ds�*��g�K���pg���
(/P'�P��\�~���W@��L����y��|p ���7��_�T ���T��3�jA}p�?�S�7�����̸�s��+z$�)
M�M~���/3K3JV5x�KnY� -���a��]5E��< .���\�<�\�Ϡ�>hާj���ցr�嗜��ٹ��S(^��ȾJ��!};(�FE{�3osG<�����鄓�i5��Kg�5`��NAX��m�4<+{䒢��;m=��8
�~de��yJоH�N��4�A(�H��?��Tڕ���̟�����HX_�+	�!C���&~��Jz�췅���l�*%PdDx��O��O�*&%�qǝ٨L������(Uy��Y
dH�����\�	[m5Ax
\_&�u=�#B��ɥ�c
������O�(�Ӡ��mq�ßwܳ�Nb�'X+�Bk-C�f�}�Ջ�%�<��:å����?���?L��;b�:��7p�nV"D~����L�E�:э���qg���|��目-2�,}�3-����4��+v��-�����G�c�w�|�{�I:��C�`K�������=���
��w�^�
�.���.��d��U�w�8�����i��v#-u5���c��ݳ��hl�m �h��4	{5;�qqIJ�裵�=�B?�r�a.ʰ�m�G�|A1wՄ�v��i���B�oa��c\������zO�J�d�i�
�1v��~b��o)�6��t�%Մ�!o .��@~na$���1��?��0��ѰK0֌9���= �"g��ʋ�MI;�X�@���N&;R�].R\H��N���K�$9����0�qD	\����Lݛ FSd��7���C$:��a#X�	���^-���)8QM�д�~�E(�u=�[̼��r��$2�f�M�z����D$�[�n�y���X~b&{�*��ޮz������K����螜�I����s��7`��
�W.���cЃ�x����w;��B}�K_��&a
uF5f��p+`��B뛉.$"����$��(��"�������R��Y��\R�GG�5�0^���'Ox��ꛎ�GJ
��	��<y�T[$}̾�t���k;���O���o8��gF� \ۡ����҈��_!`���V|9�a�Kb����vb%\����0���q�dKǕ�+3����e^��a���}CF�S!<Fa�����b�\�!x�'�E��N��r峖`oJ�Z�l���LJ�;G9�&l=:&s�PśR>�sm��;�7��x�}�����᫮�㓂	r��� ����3�նw��v��!4j�w�l�ϡ(�B��,��Q�Q����H·���1:ӯ���vX�ylUB
�dp�	�W�>m8O�s��U���eÚѲ�R��'rpٮ�얚uǙ�ϐ��_T��(�\� ��=�Đ�i3l~��C�g����H�3��3��~���Q��zѧ�N����a*RD �2� |s�U~�V}l��ByLn*+�V2��8��"��� Eo0�jN5w�ެh]��AI�mB]/�$��Z]g|[��'���^�n�a�[��Y�z�.���<��4�����zzA�����g5]�Ғ�
�X�A~�TZ {��aژ����������I��~[�<���;Rp�D���)�@�wI����^�9����a� �2a�.��7�E��q�u���g�����>����?R"©6F~!sx�?:��)��{�] R���AN'�M����X�m��Y���EeO��]�-����L����}�㊡�Q����`¡���� ��jpOx�杝(9���[��ld�E������Es�bG�	��j;��Q�vқ�MƣR�s�4��t�c��@m�����	!�r4��zcy�f��\
�Q�l�~����*��E9��᜞B^^'�[�F���4�����S��xt��'��I��gX�E�y34�6�B�Ǫ��"�vg��n���j�3i����&�y�yf�%�C��Z�p��(Hg���p�+�<t�4��#s0���Y�
����ɟm؎M	�q���nK�8�3�?���p�?kW��~��cy�=���nB]���W[5�.���4.2��'���_�ی3��쯴�u���������)%JS-ē�\b�:�y�2� )�^W\P�z0�vp�p~����j)s�L��Z���,b�z_1�2�m ����˄U���e_�^�!���@t��q���>A��3`���M��z1�3u�F�f���\��1h�I����2$��#����՗� m������|�W�Gם�6�}WV,<t>��>s�נO�9�Wh��Q�r��k���<(r���M���f��j�w	*GR�Ultٸ
�އ$X��xBu�j*@�U�^�;Q���m�M��2~`�X��cH+Ǧ�����9�7�l���/��R���i��Beܓ<��C��Q�~�4��S���6�Iͤ�|���k��d���h����Y4G���zĊ.�	��RS�ro�̬����d���Β/�>�z"g#����{	�.�iƠ��2.������Z�(P�����C���O��2V�ӶI^��c	R#@ryJ�R�	���ٙ��^c���'�0�.D�&5ZdF�\6�7
#%5����b����&�rT�ƒ�qc]�RNz�4�|!�? �����f��i�.��u��^Y���n�PZG�z����;���g�^`���ƾC�"~-u���Y���% �������6r��:�������8�Ѩ��c"��>u�P�jhVt-տľŐm3# ��3)p�ǎ��z��F�t����Yc����k~���� %Z1NE��8�4�u��]r9qC�}�ۖJ���1�����c���Q)�qI�a��/����|��v5��:�8��3�Q�Ò�N2̄�i5vZ$&[�,��t#�.��F�E������Z>��S8̲��vB;�-��j#��qܨ6�T(U�N���ڸ?M����`�"R����5d�%H6��9�$�J�wG��๡�5�(�vꡘ*�[�_DHK�MTsmmR������_N�Ԟ(Cހ��T�<|D��w�ڊ�+zT��l�u/i+�k�gY���%/�Nv�5��5�\���	d�Q�8M;N�c?iL μ<��'�&ɨ_͒�7�V�����7����~����Fo�}:���OHm�������4��d
F��3N�_���~��U=*�ן�L(Y�5��%�El	�X�j�;N��C�+G$�b���ǎZ����8�Br���i�4�I���w��=:W(��8��W�*��V�X/k^�[�M'�T�lFb�]��$�JA_	'fgF������4�(u����
�6AմJ���\FwB����dw+��nZ�<���]H�L��P	�t�S�� ��&����0��P4��)��o��
�'bs|J�K*�I��ݸ�Ժ1��UW������(x����&�����'(��ډ~K�m������΅�a��{�\�
X�iO��jW��p����M���S�}��B�c�1��+ܙ��k2�ʲ9�!�L0p�:�M0��!�c
�Ҹ�B�
��.~������F��#;�K5_b]̴e�Q��\����c��w̞N����o�!�Dީ9Z�&s��?������Np��I��H�ai�?�
��0�C=7��>�XA�"��O�݀?����^����;E���� ��P5��M{�5�4}}��2��	|�7w�j�W�=�D�S���L���^%���G~�t���8w����8����A�2�J'g"a2�c@�e��8���[�C����#3iV���H��
��b7�7_#�Դ��D|��O.��!�0[-G�*{�ND��[���B��+e�h�b�n�����ih�s�C�"I��oona%n�`�H�l=ҧ$�Hs�x��,E|�kgD�P��a���R��B`�����/��]�ޠ?��Q�q��э0���[)��~x�6���e�JI~��R���a�d�}��2����&������f�,ބ�5���+]˟��8J\��[��k���םNX��e�F�G��(}`����#�8�B���h`]���>?L~���l�BFeWB�}Wo��#ץ���~d]Uq@�6�!L�ެ�.���2j&E�Z���� ������C0v�F=�m�dKEagVmu��\AG��#|��P3���6'%�N���IE^	w�Y�eŞ�1�G�F+�8t��B#SIH���ܶ�͂%w�X�?���IV#�i�ݒn����1�,��򸉃����r�qU�Qn��jzgě�;�S�[��`�ۓ�� ,��W/���1U��y���Er��Ŕ�75�l5hkn��`M]�Y�]�*xA&���	�G��>f���H{HX�䶸0rnȤ���̭׊^�V�,��[3[c�6��M�u~\�8��^��ʚg��q銪�b�	T}U�L^��Ʉ�$cQ-N��ʩuՌ����bU&kV`�Z�0iW񥖔	W��3/���W�{�V��OD�	��:��&D�I�g.%b���
���[�E:�F.�@�s��7�`b����f��I��f��&��K�bN�o����X��aO�觀�.W�)��OeL�������� �����hEI�J����mS#L���K?7�x!&�2�:
;���~F��Dy\����|'x��X�8��E=}e���i�]BX��z�%�N��}��GrHH��?�T���$��R�wC	RGz2A���=���m�\�]c��L��B�6hHM�^������m+�v�	��n�(c�Ih���`ѭ�i��q$�A�U"E=G����{ILRE��͐�����F9�?1*�c(RI�"��wt	�G`��!�"n��R�ܪ����A���:���k�h��UV�1J�x��j��&Jbގ%�M���)�taJY���};	�[m�H :��`��Pٳ�Õ<[��]M���t�'�\5Y�����\O�%�uln�B�ӯ<~����c��F��JG7�ԧ?��*Vqh�Ma34�|oh�a�� �\�,v&u�{�k��.�Zr�%0J�*&8˸��g����3��]�cy2p�'�3�C����N��$�ܴ��L_����zT�AR��8z����RA�v�z+�
'��>H>rܙ�Z3����Z@G�T�2tݫ;�ʊ^�D���^j��.a6^���u���R+��g٣�����RB����2sJOj�yv�h1�q&�Q�5�v=s���-]�9�|�+]'�%��g�?y��<e�)ƥ:*�n�^e1PQ<j`�� vQ��/��fIvjҿ��4�xK�\���eܩ���6Fu��Ȑ-;J2�ُ[�TW��������Y�P����Kn�5�t@}o�(
���㼄 	?G�Ĵ�Rp>>ĝ�֐$Y`�.o(��`G_��������j$�3����A���&q4��	ϻE֧���<e�_y���F�p���|�/uTJ��B鶨c>-Xhj{��}(�1�V�0������i�������Q�hb�MŮ��t{J�ԉ�H<G����DA^�Ɠʮ�q�	����a.u�M�,Yt.�Ѽ1wS��gY�H$��0��<�!��(�4�k���� ab�jz�����������"*�Z�O�ĵÐ��!1'%z�]el5����\�¥aP�ݨ(4\N?@�Bi���TQz�c߈���k�(&�<����:�TW��3�;�['+�N�li�
���V�~X-�'&p�ǀY\ VX}2'�4i��E��ϳ}w����K�u8u?���|7<Z�Z�qd�@,|~z��~R�q����,
�WG:PO���v��n{�!~�<����̷�3=��hE� 7�������&�����l���!�1�`�B�{�������D� ��ʧ<��Sg���ęL&�ދ.��P*�H�t:�'ڜ�~��sD_�ȭ��,���<�E�e�y[c/�x�~�pÆb_�����gX`�����kҎ{-�B#��z�;^� ;�c�z=\�G`i�	�k��X���ӥ[��i��Q�e����8"�?.�ŭ?<�lB+K�υ�dm4���K�,�W�RZ_��_�'�X��f���F���O3ju�a2�G��2T�0W}��h��ΰr7���~8.���+O��fET����W���ǐG��&a�|]�L2�b͈#I#����+��ȐSƂ-4	j�,<�	�����Z���;\�~���m\z�y�Uhf��n��� ��l`A�!�[�aa!�o��eb6WH�c"k��G�A�N`�.Ba#N�f�GN�^m\�-(D����i6(��Q�[mG�=���
���#i%�Z=Qv�y�sŵK�J`��q,1��}+�F���	\+V�+L�`é�
�F�~�]9�c8�-|�Ӻ[�H#��7�V���|B�����3�~i�m�<��y5������d�r��m�I���C��C��CMӕ�^��g��і!=�jqy2�VQ�Y��+Ĺ�ܩ��r�c�b:�J�sQ��?$2�Z-��zy|�x-u��~WT��6�uݠ���h����M4��F�~u� ���E�D>M.���W
�8�yt9\�K?Z?��d���~o�K��~�s�����q4��f,m���skjMd����iq�,�ɀ�ު]�=S����v�Fv���K��Y�u�R�&湞V�+n|�&1��y��Y��:��jt�u�#	�5]�����if���t�] �#����z�o,@��1L�C�2V��r��=4��`
�j��e���q�\�2�rj�N6�p"�v=y��p �.H�]���<Q��H���B���x���3�^gP�|W����P=�֞�l��cOZ.d�
#�2�[P��&r	����� �:�_B�ơ�v�L�q�
R|���A[�~
g�F#��MqD�y�����S��F=��ۚM/�.S���f�V�.�o˗8�U����dLch܎K�<��/�z��M�C�}lɴ|h�f91��EpW������ˆtʖNۊ����\1<.Q�R=5��[D-?X���2:G������K{J�+���i�^���U�̣�9�Pb�"Un%O�=M��8_�a���o�A�MT��m;���A=���0:��r9m������`d�Q����v�����]��VRbC���Q������oe���*2�s�VL@�����/��#E�y����9����[%���-:q$�炱0����^�P�7S�^��@�1*s���j �q^c�2��c�(��J�y��s��[g|�
�Q���A��)j4�@��^/�,笭�]8[�b9���䂁fUep7J3���O�R�c^���SY<�j�	�J�n ��Lݔe{�� �Į7�}�q�{Pm�v����2V�T�4�pF�����C62��`�e�j+"ܻ��;��}<F���v"Xj�������5z
l�/凐� ���m{)�2%^�r`�R��X5UJҲq�Z���<��,��I�/�+8#ZyZ�p�j�Q=o�/*OF���Sq�}w/�ycJ^���!�ևŰ���[ 6�H��)H��8L�ŭ���L�$\��x����Ԭ ����p�Q�U��R޼��zpq��8��e�wm��:O���AH�X��9��.;f0C��9)f�"d�N�砱�ڸ��ٹ��e��/<I/4�^�����bwɋ�)�/�u�,N(/�|�#�.��5�u ȴ�rؕ��Ks��Eɔ�[�}��oӳ����<�/��:�>w������ۑ4��1Q
���o�S�G&�.�պ�� g"v���Y	��
�5�&���������J���0�su'n-�傱C�^I�$$`��l�ӵ�cN%�5#���ˇ�$�U��8�(�� �}F����b�����g�{Yh����?�c�	�P�}�my��|sO\U�i������JD9O��b\�"
�Ȁ\ ]�?j�4'k"����F�QBgF�bn�3�d'<`�C'M�~0y�TD��X������'�Գ���x��#����� S��f�s�`�2�����dM${n`&o
}Ǎ��"H���ҫ(�"��z��X��-"&$m�:׮d.~7�Q;���tѳ�i�hOqE�n�aS.CmQ6�Q��8z���f�����#5�cvñP���hj�A��&�X/x���;��9�� �G1��0xX=�߯N�V�mN�;.V�/� 5�5	� ��=o2�8�|^N%і�{N�&��&j�����#�LI�c��_���������1��8S��oic��޴���W@���)��ʘr���j�m���d�#5��࿛���p���绐dd&T��@�D�䪒�ф|}/�;XGT�6uh�Ũ�2f��P]����O-ϖ�/�$AJ ��?
���C�w0KѾ�pC���!
�O�c7��{��ޗ$�߱���N�e�e�����:�q��������8�JR���-��BbZ�����Ew�4v����l.]���`I��:J'��1�`�k��F����Ç�P����/�e_�ZcW��������ۗgm��k>>M�
����BN*=�8&F �Mc�I�*�=�;�3_1�QՐ�ϐ�Ƴ+�M���X��}�3'���U�쟴C�oD^-��(3��̺Jg��0�o���_�� ]�;o%��t�y��������u=��	nE�i�Zl�i*���73tt)nVX2��y�˛xyG�Ъ���94%>r����6B�c��N���4�!�NwP�TR�~�!���u�].I �g!H��b��B�X��o\��X]��#�_���b|�����E��EO�%�'�P���ς}E�*��m�s�3usp�����*(���P��&��G����`��;��! ���Ԡ�:������du�T�}��w�
�̘����I��jk�+3;=�n7�[�I��e�̰�J� �g�