��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2i�>�|���B��,<��\ ��W�~��O�?��K��<$џ_�!�ʙ�E�?vo�7O����#�^N3�Ny���,��ț��WV�8BRc�9�!k�������J����	u�<��%�r�
|�}��5���ϱ�y03A�4UW[�^��מ�!�3߹�-�3gP�ǎѝ��T����� E�}�}i܋�>
;ȑ�Cu=��H��Ih�VB.���ls��~��G����P�� g�[��1U�t9��k`�vI2�����+�1f�!���b��3�&!_�}�aT���.N��%��BP���i�%� �����1�G'���.��M:�e����&��i��">C�T�����B�\�v#T�[3b�F����A�Ѵ�n��t)W�Ql�|�T�N9�Q	 �/޼~�<�2Ll��wv��n�i�&x`�M�_W[DT�i���~�3T~u`�#�ᆳ�yy�h��f�y�E�������Z�@Ə3�*l}��n�G�t��ku'4���3��ޘ�+��En7'<����i!�����öq��G)�������:	���/>�,n���eo]%�~�����$���g\��>4��ї��Ƶ�-�J�'�v��Y�x[a��qG���oI�d�⇏��ݠ-[�����(�'bn"I�W�ćh��UC�eп�,='mv�*�a��Fh� ���=��ݎ��
��N��׾��ᦥ`}$Ӻ�ׇp����u�N?5�x�� �n\л?����o���}0�mM�Ti�qA�,�����_��?R��O�~&�Ɓ�y	H�b�2�g7�ѧ)0Y��mת�4	��6���9���,�._�+�N���j�j<��o;�ޕ��z|�9{o���+[a�l֊f�@ź�7����NO|��F[4�����6j�zs��/��/��{����Q>K��c�q�W1�y�}���}����g?�)�?����LX,�S�5?���'���xQ��X|y��Y���*�b��y~�"�����˙�*�Pi\���_��벗ԧ\]~]�7�nF��N�+�\�Q�۞zҔS���8��۴Ҝ~W�h�i�>��vWa�R�-�Q
ip��j�a�J
hô;<����J���:���lXa�7��9 �#�IRt�GB�R�=� 8�RۀFb�ͬ)���ߏ���s�ؖ;R���q_���K{p1��*�v6ao���G�͆�a��'6i�z��.|�=�B"5���.�B<J������n��uO��d@.S�����k`�8�?/,�����jl�U�H٣��M��U����s���")S���q�WU�	I{1�	�l~Mv�j8�7���J��h���Ǌ������Ն��� �W��/�w�4Fs�i�ۮ�4W���d&벃���X������)F�r����r�Y2ͳ�I�$t�"[�	o���q�� �P�bX�,ǂ�[�-
W�[n[�&D�T�1�Dl�bZo�poԥ�����Z"�q��Ѷ�g(��4��	�!U*�y���v�L{�Ú�}mF�����}b=/��gi��Kh�/�g�s�ƈa]ͩ.�GJ@��eT㕌���A��0�o��	���{���~����&\�/��!�഻\��#V6�f���I�#G�� �!�xvi���$m6��HE����qh?Ű!*�N����f���`�A�6����[�b<����*EQ}t(�N���J�ĸo���W���g(r\�������+�v�~��x�Z�Hl<8�:��7i�ɑ�ڷ�C��~p2�9V�/|cp��|H�iK���^Ή��j�]�P���d���*�f�2?�G�����(���g�Ak��W[�x��e���6f&��"��ѣU�,`+��"C*��Q��0y}�f'#����ce-�.��ǳ�к_���B��\�đ-����}�!��G�f<X������,IU�� -m��Z����%GCB .'cqi|��a������+z2.�H�� I�tIR�������C�8Ѐ��<"�{�@Hg~�TJ��=��-�üh�Ǻ��w��հg���	l
�R�빚r��"��`���3��5G�ۣ��O�k�#@Tw��O����H��6p��<��ityeR�O��,�T�`p�[0����W�$�=���E�^Sk$1�\��!�-f��G=��ݻ��ʰړeg̠ߥ����n��9�I�U�IzTsB+�e~���o�T�*O)�/o�:J����l�b��I�}�U���,�]Vk��������s����Ka]*�nᄹ9�)�rL�#�	�h�5���j�|;8i��BR$��MZ���#���[�i5|�x	���������M^�l5��+�_)+m�=�&X��ĹZ��^�c3JW&d�h�Aߚo�E4���,"��$��f�"���ds��jB��Eb�?T(�"����8��{y>��hA����hY����U�on$��`����b��м��%VT�L�yqm�Z� ���`�F��3Ih8�o�$��u��������n�S�L/��U'|`���#�&�25��U|o���=hf@ClpU�g����rЛ��!L�"�p�E/`��Gטx)`��)  �TB��ݦ�v_�^?e7��"�d5�uJ=	S"j:ǟ�<�IZ�)\a='���8T�Zy����2p���4����>qZJ����s0r�燂.�6���%����Q7e�̞��O>�I�ҘC��=!��\[�g�ۭ#���#W�|����s�;�