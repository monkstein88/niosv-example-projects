// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
d6SGwy8k4NkM0Ww2EmFFhD45lR8qsofk45hrF0Oj5iBJsZEYLfb3Cia8zxe0PFcpplqwAchWuvoF
82TY2Ognr1LvodepbUVwXuQunea93+UEpPU2EdNVDOq1gHiV5RH02n2K49XFhxI0OXNPXBwfuO7U
jqlWvdr1il8basVGPkqJVCUWjAB2F07MgR+26w3wZ2ZFT0oOaHQbaweKIjRPQDtSGGobUM0Lz5lo
X9iF3uTw3yt0jOg1zF2a2N8+TL3eZWmxcAKy6w157UDfCw7Q6c0ZyQIw4hWkhbjR45OUT8aomWq0
IPhBoWhF0jjNqW6m4sVgKNObSM2MIZD5un9XSQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6176)
egINMHHaHPhLrBWDiilLe0rL1+ate7ACU5nAVahHsnTmbJtElmnffdRvRFg18wBGqyxItdho6l5C
hywLp60+85uY9EhhxMyB0dEBIJHUgFGvHrtnAS4EYNvubkKIzBF5p1vxbDvXeXeyodWvkfDox9P3
/E9FYku3foruml3V5onc8nopBNphjzZttG8azFhTw9c5ETFMmvBZ+KL8yw3/SoYxm4kNG6cy/jMM
X04Tl3S+bJb8rnGPO8mrI5fePaCTR4uRUevXSN7xgTFowlAlAgEM3ufVNUL5F3Q1ObphL/n7Wa5k
43BZeGVq8P7BR8zltBx5A6gTvCnNVkwvZOg4Vyq2z+QVcipkDS6Pv4RZNAcYQ58AtTO/Jy5y2HzM
dZjeGHQ4NjHrl2bohIb0Fe8Q+kClarnkePsP3GilPCHxcPm+VKKcpBUK4O4NfafzEakCpZD8V+9B
NDAx+/daw0H9QyR4CLHYKZwQrd/xWeY0lsjEr0C6tG0Jq0TXdNbQWwQKjXNvo+HWUxjtKfIg6Rxj
OssgDkgY3+1fT2fQ5OvDf4H0sL2c6rsDBOsMRtISOtCW+EmIR5m9Nvb/7URJVF0iOhxsb/mpbkuS
TO7psChsXGsewrb3Aw9D6BIH4bitWm0MN4dKTS8D+Cn6YQPEb5lEJBMxwCj2DXmJjmsfjMkfRvT0
GpeiXk6xYFDa7iJ6O2C9omEOEYAtI1W8XDzrXGShpnhLuTB5Pi8ZF2JC3Ndms3dFMZ59cVAPuXjz
J8vT5n8I/21C9e3INSek3QqECpy2HeKb+24Z0eP6zpA2B3jXqpmrrgTX3fKFwA8MHSsF605zvZOL
0K9KDuFy2WWCeomvog5LCO2O7s/FBn9dhfxU6Z3MLtaRUaCBOJHaeeg1aXPd0l41BBjm4n6N76Lv
3hj4Uojr5ZFV5HYjubXKvwGEg5n0NFR4riCnvictcNHX0bDfZLucmusvJwviVWhq68uXGHx/yYIJ
oNfidSgykfGTJ1wVPapSRflpC5o3xwgRSBt/B88UOXquoXVV6a2xikgnFcRwlwsfqNnwhfOXS+yE
aZieAHyanZe9RhR5lpZXbasRfDK1JDQfeYf/6G8yqk/tV3xYaUVctZzbuQVW7ktmJhgzrbwa+y9j
KZXRhcCYJzzjKkcwzSwuUZw1tV30PqawUiHjeQYfxL/fNxMgpHmtBI0WDmciy1Zxfv18F+I2WFq9
kEq0MTkdQPp8mDF31f7WXeMhXNQtj1kWxS54Fl5reL5tj8MHBBORZxvVgrmSe7zopy6eWzipNcp7
5Rn6F44OMUNBAilrljwxbsgrDO4A8UzJcRepq1V80HNKhP1iUM7IZVBpkJjkYC0RjQPtKUSl/QJu
0Apql9mGIpm7KcYhaKGykItE3ZyF6pd1szCNohE8JFHnOAmnETcWzWZFthQRPMS9rRILnpJ7zssF
C+r8fI2JRfA2A+Ule4s7XDsOeRT3pZK0i0b3LKcCFbscX53DSsANwEU5u6m3OYnsMyY/y9rNJzit
VHmJGXS9Bt/DUDO/XA7ruHV556CpBa3GfYWD8DjbnnLaYCU4e2PiwqvOQI1IRb1zRKWOs3nQrh8P
BNxVEPiHi159o5VkF3p3oZqaS2nd0BKb/ay68cDDi/iXG0/wxRBYlBxH5nPN0GsSAOACMSelyn/P
6UFWDHfNETMtIfW6JYdep+IyO9nYroIn5SBK++/FrqcQdCKI14zWlOKe34WY5AygLyGw1Sm1jho8
O2Y2Ch7Rfks4PwoO+5XEroOUbQHt1wzLse4fpjIQH3B1zLa7JUA99+5aHG81jkTiT8yJ71eDmOn3
MngsjHmpnJeXhhki7fM9iCxt4RcLs9yOYWUra59ynyFx975sKDpC2BZqpBpqM6keruGXxfb18Kb/
3+dP7kAp0QLYhjwahzZ+dQyBdtiU9jA5m8qQT6BczLEaxsq3hz6QdiIfGsFOzSp1cYca8E4BGVHh
Vd8XaCR5OEEpfCT+pIhxK2sCbZB9TC8OJ18h3Tro+jfhEwivyFIk22KkWUqYUPExCTURsAmdTmAK
xJqEZnC9X5wHsbsObX43WFwAcszaMsz6U+AdZmTSCthlnWhdOzolRfizClhB5mGjlenZpRanOanV
2oQ72FpDeyqOFH1FqYNlCZDJka1gj5flZquJdp5Q+WR1uM4OgfV/Tdoe4AfSvXYbL+tL9jz6efLV
mzXT2Z/kO+ngiNcNsEOhXwFv2Uam2yiu8/CN82POtJq+bWEAaN5px05NKHgKEWBTRTsSm2Cd45vu
CQu8vA3RlZE/FsRq7ku6Ixds/1yiTFIGm8hwdFiNfJKpbgPF4bn1eEWKDLHziC5/OXqjoNb+W4oA
Bxj8TsszEH4BCFEbtrE+t//P3JKjUdgN8VjGl7YVpytfbLJ7FmJv+Q33qnx0fnFc7FQAbcjS6+ee
GKL4WLrFtBkUqVdfHGkPfMiIrTZW3KJ+kXfEEJ3qG85IYqrWMU9J0qUmv0beigVp6B6I9le9yofd
o327vL7evDwkd2xEDkcZVkVDljR9sjs9x8Yd0exjnUmYp0LVhhOMrqgHQ43iBq+jOGbwZoIahmif
rOJJ6nsK90kbzaxL++ojqL8Q9z4113qyAmC5TzdN6qGXmDyFU9txdgCnnRqUu9immErgebm0sO+r
XtDYebOXBxy20Gfn2pzSV7n+TCuOqAg/beBDQ449Akwhc/n7D95mI9nq6YPIT5CNfg8+fsM8Kiza
j1EP+iFvSc5/T/cGb6SXVb7vbsQKRvZfSRuWUs1elKsWapvV/hDqYVgoxuvQR9wlQhh8ltBq28cl
Rlpe8AlmC/urZXyxATfnMaH2WOrYmBvGtnWtJJvKeq5zpgX2jJiTjekBcu3RJbbdc2ZqK0lKQVF8
olGTbHO5N2fd1aH+X6CF2kvHJQyTH9M/vGAttTM0x4Bl7VqM2bKVLTtvN45OOP5QvR+7RAQM5Mbu
WVAvx32HNy13cgRzLuBoIpItoGtSizQP6WAZGMEcfRBVEq2iILgj6tK4fHevn55Z9JEd5237+QeA
cViEbrQX8qaAAEyDN6/+tOnfCmty6sgi+tuuddrVlhopS5/pbYibJRMbbY1AX/gEZHWLGCK6Blgg
UftmtAFgrjKfuJQpjqtoHI7VrAjajeH01tfBnkAxjHPCZLHllt0OTAZJpsA73bRJuZ77R7o0+ndo
IIdX+9yYMM3ZKDBguNX5HH/WsprpG1cO+j8o2v/F6pmB96tuh7uMNEYA5k2cKbHA+tJnZw4Fw0YX
3SjhZxI6ICC6RU6qCFh77HI3dLyjNVRO/S7ebBXySs/Pg3ZwaAKTec22dcUYgVeviPMnYJ5c7O/c
gdY21tPHqimpdEs8AAK/o3x/E5U0Tw61c+X+CwZWHpCQtiNeeVbR+h1d3im0ME58TNu1uj7isREj
zqd2ky13DmagT0l/h+QoGB+BzNb0NbAkir24pojtw2HXzYOKdJCNK6wDt/Qx8t/DqqrwWNeyIgPu
lFdp0iFaTz8Jmplq2AY9QVRZ2xq+ei2xcwt74IHXV6TDpupvZpvJIg/9lNelL3HnpLwE1jEMiMUC
ZwWewoFzHLP0kZWLLejNA9G+/yxU525AihiA0SY9c2yNjCp6vhqyFTfDbro1aktqDXD46zch7c5Z
G917sHcnK42UNvGPQmmhyLJQI7g4P6Fz/EaUf0K9x+3gDbGuVYl+injzsKL9/u6syNZC3auhODnQ
aryi9eKheVLqH4SG/xh0fzCPjRXJ35FhtxZ1PgohjXe5mbIwursGqOarLe+QpYFjY+OEDgx2sYyP
KLDUvgoRHvTiw7wVUPcby4YQqeCHohNQEaoI6iNARIXdunhPQCCfBDlzMK5ZHUv41M+XSlDAbwrP
8Mna93pJCX4BWmciNanSR4U6s/msybNLGOcNqF/EEXdZWo4Ss5FJdEMh4/UU4HJT6skPl3ciGoiG
K2dfzDMX15I0DpkwbkarjFF4EghuywIdqR4TEI1x2zsbGMNglq3HNrxRErNj2GhsnzReefskROrp
Mc26LyfQ+hdcxiW6e+V8L4Avww8mTVEfc8m+FDU2x6Wqgf8rOrAiwaHvo7NmBPqaaHntDcUxs+iZ
oLb5b339WbOE9w2ccbf4fsU99UNMNk3jzlp17+hB/4GQHzYmsoBKKbayelsBSJRT36+hIcFA0lKk
s3B97hdhh/tkhMcSnoEmKoa18sGGL4O7UR8M0mLG5et1TiQ8IX+f048vXX1r4bHs97OCgP4eSGwv
ecP7ItdjfcG2oO5+Q0wfZ8FK2w3MFAAemBtMHXpV/CTdGrWMAQb81kU+WzZF7/dnTdkbXxTOgHl0
ebYuV5hvLFkqHjj0GXfe9TKWdk5Oyh8uS6HLEDC6IMbUnmt7qKTU6IDZG4wkvSF/ZR2n4sHgIZto
Tp4yqEwgXuUFNjSl55Fb7dLFQ172OND3bS82Im9aGsYi7UvcdPncUetzg5344XeA1qDAQAEDsDKp
NNOKYmulGUNp0HDOnswDiJzkP21WW1orFMtETvhTN4GMWaAQu6ZYf+1R0goDE0AFLKDsUwa3KOCc
momUPlHMB6dLNUY15U4aBOVdQZPepz+Vmxgf3G3yliqi3Pn8bRQ21DKCZtezmmGkWgzgsyjtdPVr
hLUeiHIdQKvm5aWwJVZ8nxVTlnOvx0DBJRC9VxuCFK4/OVyEgJ6BMuTjFJfTLMIv+hrgNkN9htAT
2mwJEeaVNwJj/Gn660r55+uELtNv3X39IppZO7CzrVp9RgAxJuxRjK9OCkcSlW1P/CtEZC7a2Huu
W57JH6rzosdzkF5q2WZK4hoyecqwlJylX0Zlv1sTjGu5ay4El+XwhHwYSqYWx1TuXz1mLju7BnBB
rq8tBk3ixrr+dx3BHo69UAZAYkcglClvCLu3ozxSa7Zo7J5VKBjRfW0DnS6zXRMsR0BHvkDkkxL0
50bqWrS9WF3l3tEwJxqGzeqvRPpmGpudvsr0zwTP7dFaA3JlJuGhefM5Dv1t2f9SaViP2GwofL0M
OJJlZ/wBBnBoOvOW4H4Q/c4/uYOBYzka3AaSAUx4DYQg3N0vPl7o2WeiRR9WSOBvjnNIL8DpYHwJ
dAyKUhxokKtxuh8qMutXajWp3hpBt+yacT8Nc1bZ5db8TZGt/bf/Xx64PmkHhvzGxvTxuQ2Mdmzc
5lMrZ2YqSFPTXNpbMxWx3funQrpvYfaVByLrWzHRECfnQhZrMgmy2Vt4lLRBG5+zqgQff8lzDniw
O8EZ9WZVfQ+3bSs8y1aY9yi5Pi6q+WC4s3PnAmyBpCmZccdenR7K6ei7/lFmuX37BlDySggxPhbk
C/ymF30bVF2hFDBRIcHZ4X9cbZ7byHWb1RjpwLSwl51uLZBBwwB3Dcens1/z7XoOWCwrVyeRJe9W
JnNt2xEDIeFJ8keFQaq+b13VP/Eu11iAPr7e+JTAZYndEPcWwZlsqFE/L7QVVDXCFoJqbTe3K9Ci
lxNy72CEDX5JKmG/iPVh1Xbx0kaCS3emuh3I21RMYGz8L3Ts6BLFIHxJF4fRj4ZRF6vbEh+D5RlZ
ZIRKzAT0XaymycC18fh8PhMy6U1dBuiJWTY4o2c/5msIHNW4X9XvRX88GlJpkwTQNJllzJeFBmuF
ycBShq45efEsctKaUR+K8ab/ciA31xA1UM+FED8ysy73jY6VGMt2FjsqIDP+i0y0xjoz4WDh/vPR
BweI/ZLs+mrTWVmpRvzz9wZMCYGyTI3GcudwVMVf7WcuSMt313pD5Ow2dNOWgpEBsokxLAJ1n6wO
MDl6xRhswz1cLyuZu/Ur8/ipQ81uqy4cW4874cEuUkRdDxyPzThO4KduwftJZqroJ/1J5nQbKeVE
FSGZBGuHScPKYYjVUKKCXWYb8cz1si7U3V+5AHYKM1LBUvBXW4C/iXBnrdHtvW4VXsIGBJTFHd1W
H4uJP18KcyX71bCsuRwvC+6hH/jpJHQ8ES5YtHMjWetDb2guM0nzc2I48LZ4zzKDuWuU15OUcxcl
8ck+S+1yR95+eeAtn/eMGeL2gLdvONp0WewpV85RobIzJnWhQ8lGpsfDwHePv4oI3BF3tSXHvzoh
T0W1ID6oC94QeZr3ZfPzIlvSt2Qw5GUV/kVa4O2F7ekBLHH7vk4ku8Sene1qBRNVnKCk+q2czeVZ
LyGOyDQQS7kg4K257Z6oxg+VzNYjyBwIQsm6dQjuixekkxt8nFFKosPiqExMw+a8Dix49/rzRCnG
CLo8d9TG9Mo9Mh4lLVSNrM2uW1fIeu0eBn9sT4GPzqhhdLr7TYSdWiEKxCiGCIVQdAliFek/q5wf
v4QljYCwUqymanwr904NaeYnf0Mimq2UMDElaGmePQLTmSlNWzOoNp0E/tIwlsvte19ir5MsdsI7
6VwwO55a1gbNT/DZhjX1dbn+witOfStyCzN0Z7QZbQkBGoQ/knqEExgrMQln6QtCnq9vuT8oh4A0
CkP3cCUNPBpbQFnbvBFNjUGAbNIFG3MtyRCtI6jK8RDaAxX5IPNElyOSiK5eJUvdW3zgesIXbL1n
TCrlhRe4VnSv4GmbBc82BjxNEb/zI/H80SiODtvhjK7KxhhCU2rdnvL5O+wxkj+M5ZMsBUGUCDVn
HmG/hXTecxWJCIL1kqwjcFAdGi/TibpFKfUhDK1ZWTNgF1qLoP7h6W8d+Uffk34JO62U652SjcEL
LUa7tTnDEm1AdudzKH+HqcJaKJDAn8J2tUpyXmW1xaFXPO3ZqyicxKWXGUDtHFq38solwF3wiCk5
Y42c4093nU8nsPn76+wvTlHEb2Du88RdaqVt58Tm22jR2ILL1fXIUXpEvlfpd3YfvMafNp+lUF+u
ICg8BM1Hdkxka5LMtgtpVq3G+AYBUCgiw5EPKBlpDikZvEh6lPLjvMld/29tG5cQm4UA1FdBR3ze
Au2+cYRFQtdE4FHBBU71IfA7an3nRxhIL8TGMHGcRYI6DJYV8zEAo7EoAbDcME/G6eEz/vkl8X0e
ForplyHJ2vx2IcCjTu7sYxgHtv+cJUSRrOKobsg3t1joSehrhegvTSBeiN96vo2ACGyUld4/t5q7
F/y6xZBe2gcIIYcrZMFUq9bwTuikfIJg2k6jmlxPssJPIQCCSnpu63+rpf8525O0DnqpiVfmTLJB
C/z5M3njxBhdBruVEHGRdeDCr2HqvEMXosfs44R6s5G38WgqWj9EM3sLeXrKQOMYrZx1dUSdOmJR
7AGpBM2JI4UbIhB1CIIdV34cqcszVwRrZSUFkOwQ6j8y8YetJQcpp3OWWglvTW1cMN1OB8nwLoUC
HH4mplORtLm9FQmojMftK6xKJVuxYW+Mm5E+tLCoYym2/TqR8+CbX/x/c7HldXOXZ5rN6iIxFUGS
jJv+hQY67BS208P+fJzAjSGaULplsaU3wIrl3HJ97VTpcTwG7nCHtpL07JFH2ByRJAxUw/DyhlgW
Kj6QbPRTsdsVtNKR2eGQvwtbsMjtK0g7iBbn9Nw0dFTL3YkVPM30wKh7aZCL7f6sH/ny2A6JMwtJ
hYzLlFEuhVCbZQH+ZDDFhBBLF5/kPyzL1BiNdrk8s3osI42JhBuno2jmmA+pe6GRxSnA2VS9URYz
BxsNSadzdprtsnz5eVgxoxmICnnhpoZ4gdtHb0cZt7SBxrb5WfNDA2Ui4VO6wIEo8/gZCRZwOFTy
fWRigfpT9jDUr7OLZyJyEZg1DW/tgsoyjB2kk+CJnxklkVrFyeN0ywnaxEmUlrEfyoIaIKug+mV4
sEYPtrPRtuCV4xsQ5kehyaTriYI5tHRYKOtFnqk0SjYHj0vmILC0CTgUF2xmltzPCLXjlLm4TBnu
VOUS0DvU01JOZ2CItHWtaBgy7keR7AEhR0BXPRflS968CfmXD0/+IuIqej+cgYFB+ruJz8W7kVAL
04XmKV/ewIo9C96LKdIMBX5EXIl8ZdzGygPj4ZQ4Amf7VE0Clooet6v2UkX1a2i8iu7iw5QwUelS
4CW7KtROoP0aIUWzauVpptu/N40tz96OqXmKwn21yZtiFJZNphsi7760+yPBV7OOUiQTfpYJ+T7k
sheSkcHGww9Y3OC7FLqYotMypTH4Mnn2RyQIHjiA0AJVsOTADXYkeUvwfvghvOe4c9LmnetcQVtR
1HoeIlE5vQKk1vA+0BdDAo44PTAeByv/GGmKPqJVdbbeyQzkyZDMTOOe+lxNCw1puRFS2pG6klIP
GYSPHfCf38k4fUZK06bzHNvI/lo=
`pragma protect end_protected
