// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rVQ4rpYq+KphbrZDqGwhpT8uELjF/f6ocGXi2/9Oqx1vgbbz+UqMxCTPB5H1T3LupYU6hwVidRL1
vdqQSyGaNb79GXaYALT2wSyHB79GeCx6ANrc1fs75khjpqMCMWeTNclll2QSqURKCB2rnkD1A43F
CF97u/ahNhunzrnJylyN6dXLDFF2khQUjiMPONGFMj+BO9yl9QdEvmkcGh4Xkb0nHT3GfD/KfL67
44T4jSCvwPP2KLBDwDiLzDhhfrvLQBooGsfYcrO+TIYuouYBVPSXosaCVGIl9n1IZ3kA/5TeMNqY
0vmg7GurQENYOHu6I4PFo5n/T42RyjT+lbDECw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10080)
nWpS7fD1sMQAqSIc3V8oyO1EJKNIWprVWTHs8RI7v3Bs9oOW1iOUfe2UYKDnnk9CD+D1vFWZB+5Y
gTW7/HLm1ewTcuqFRmj1khxJKOao3PueX8XRh1brBjeS+bhhQpAgd/GHDdZpVghFGU4sUmMpzeRM
D2lZ9t3KrXle9yUAqTJvmjeaFv3SDmymvb4WeqHAmakh60by5bsDkS210LF3rZCqaHPFRfFn7xwD
0WZzJExwvM7fCT7irksbzDFp+B6fGS4IuRYWhMIozN03lSUtRys++X7DmNBvz6gQ6CA4P2bdL+Fd
TRCLOtvI32WC6MOPZG0er86lvCpdVNGYQGq+zL6zJi5fOj8yXQ+oHyxvAlgmYRZfyirsoCpqYupZ
m16cgw5CAcks0dK2/oPs7sJJrFJdjcFjDjaHueV+s5MyQns+QHX2dtZVP2KWnCcyvzyfUnwB0xPa
mgsOP1mekssMpwCguWadCZx6vGFusoK7uyBstGOR19l+DL4TA83GMgDiO7owNu1VAxjhhLmvQdK/
6Hrz1FGFXnBLNg6cN+XDfP16m0wXy2j3I8fN6JtUnyRgFmfoj/NTgufK7j41rLUsng+ezqkkHxqH
v7WeEha+BUusKOx+GVpwDdewHMZvPAdvw3TNMDhwZGZuERpS/KYd8XUrW2Px0zLfiJ4RF9s58563
LQvtPIQQZJmE1W386dgTvnQuImylb1WO01edM22VSTcyEZBeJqu9llj2fsY9wsxdcOt9rbZK1aQJ
yza6qtkUwR3m4cZZiNmN4Vohe1ysSOtVDb2E4CoDeI0AoGl6kxvm0r12IfcMaGmWVG+GulWZyELC
sV4yddCJeGorw+26VlW+TamijviK9Pb+fgNxWSd78JyWh+YWp4ADzyC/jvtGvHad3qagn/malbZS
+xxDLn8h4sVqRipTYcBnovs/lQ/xWIXOj7boGTdGAVhQwkAj8ObB/roIY8OJUSR5VGcNX7hyuDFW
bJETbVaRWUWIKlcIp1w7j1JWUqZe8LfaGjjLGKLQlC0IkLY6oY7RY6Jh7yMfIMZZseNp52lL5z5T
FNORi0rKJGUlyuHyyW5MvR+xro4EugK8KrMmYJsYrqbZHkFgRNEEqqV0lTnhzYvS4mCBbb+DOm1p
3dbhJwIuuvr/X27i9d7yzhmh5G29P8C74l8U0iugvCuGGpKXIuN0Nzp7xe3aYbx6mu4tFObs7ZCm
Yt0T9jQLGadTaqzpmcAsOVzt42drEnPawYOLn30Gu9ENh5LiQTfQyjMnS+2sI9zGbQOuPrXs3F3V
TERnQJbuM9S2g2/rTC5OHw2xqJT83EorlVSYt68i9rwkjazg1bU9Yw79dJP24aPkvAznfqUPgbGv
blg3dLtDaHBoTMO7w76iuwWMnBZHC5jLHVnJ/Luj+9783AREqG7gnl8k6Pwl1cJpAccUvGHhurB4
qI2e2GFmGlNiSgEAq0ofXDYuK6rSlz15nwSNpYCxPlBZIn4DmBk1QfgYdvGzk6bCwGjLSlpqrLcE
73OPHEtkTLxhUUUviXmnp6XmR5jFolMqrkZVmc5ju9ggsT3B1LGQVT63ogfi+ilQkjawpjEibBVX
x5adzg4Zd6nnbnVPOJswbZVv0B9MsbQ7Y79CPenvvWLUWvyk05ZyEhTKFImgRiiqP/BUlgCfcdGT
4OrfyTNHQJ6VMVllFukffHwE1KWIa5MTGqLRmuedq/0UthebFBSlV6S/4dAZ7fY55NJPkhzEYvMu
LnIGnP+UWZPyE3P+UL6DYDtdG8LS+VLBMayvdW2Fj79Zj0kx9HTz1b5UUy7IPso3WR7MLYK9qbbH
isd8opbrgMs8gijjIG+UCAkQrFGpsOOjInZs+itU9+AwwNyYj6cYAGFaBHBzWtuY56X1lZ021qbU
K5DZA/uyeHWL9GEpmFYhHVbGEKW75kTVLVdcI2EOyQS0KrGfy7+l9NxFJkIMCHFhG/eTice0uuRN
z3p9Y2NnXAss8dLKxq6vbrTMIPPWOs/vGd13t9BTBEdIQ+igigbISJRjGuBvO8sRexkoVQtGv2BT
4b+tihja1u9qOxSb9FeGzM1DGs5/VRSfXjlLGV/8RYvlgflQy318o9sm39yf2MZTCG6SYvjKOzof
oAvVgGNoZ8vMHdMpCeoWzPxAh/5BC6WV3f8EBTfd180v0Rs98Kqt3OtBAWRrHHhZjvrm/VUiJx22
Pm7GNkJOmNBqv9IRgGjVyoHfnm1LdvyOrczgRx5GN+PMK0wFqA+1De52qq6bwGRGL6I02oJcNsnl
oTo+EX2HuD3LgHvRCNlmO3VLpCECppWTAbbiqz/5wu+5hou+95akIUubmq4sB+qIuV4kdlQkT+Lq
wKb/cau4NzrdXR+tlz8z8UJOWHaLvbNSOcFTEbFG6/YrfBqe3rvuX+H0gxxiw4UWRqL+WaPEzuTM
2ycfhywlDZcNu0NqfJrTmuMvDMIUFjan9yerGqXMDVhiHj0JOz8xveAWUT2MUe1sbFtFloe953Mv
z/o3rQGt02KV82HeKYN3cwp3cl2zg2MNtrITDTdrORXA8lWRU0USA9ByfwLW+BUdDN0f5geXpujJ
0j7Isq3OWh2yImvoz9gZJxFNmUddg4XLejKWjg9CuLU1UNYdRXZSXN8vvHBK5O0NirRIW5v7X3Bo
odjieEWHx1LOaNLPrxo254VlJpCCEtTbSzb7NtCuwAXQ/ZBTsvuvjXaNQ/oYJ0i1oqTB3fOZc4Tg
JJCt41jX13fwlo8x7r+Zrax7Ot0IgOwzWGTNAteWI8Ed2+vARXOwl7SkK2DOPP3qs09k4ja17H2I
Wv5v75SeSXNRk+Yt4yN/JlX8/3B49NIpkOFoDu8hy+1uZ2R5nib5Jbh/HCUdV1bLZ8UJBQG7C2nA
Ssj+wIgBc2VgpFn2WGdYC14AJPNYnQlR9Jq4hUtB9lKZuf7TXxTIjtT2fjY00wkGOD442tIj5+k5
1g4uphPhLfDcquTS2Mk5cxyX8gsrMZvWj94WQSNIh8IO3b/UvnpMdLl7JlW+wP0dhDZ9pgi/iCmK
sY9zE6luJNbeD2POp0HjrqFu76wI92jjPpP8Wuj7OpOnu0pOXN67KCSiiDsAEVai2qX651d3rrZ8
v6VTlZEfC5pnhq1M25sTmIT8yqeduMPQLbuw2WF4w8HGl9z+Z/VLRebVDf0YSJlZZk7qLd9q3EcB
cn5thkkKDkSe6/xbvilCnNQ0MUrq67qyhwRDqZdPa39VTZMg+0raqB76bPRRcXGxl7IAEFeXyVZ8
Kb/RBWo7/Ikeo2qZeNwWp0qyPBI4OKtz9zfwosyXiP11ffiLYCT9t0YHDEHXrfxJ/3mtWADUhZ/j
fc7nHmAiXySF2SjPzdIrbEYfON0P6sOUHkoV2y8hf536py4oHo613ra194BdXgeiqjB8PKOSdBFw
UtUgjYWU4ysfYmDIcQ+8zv+2Cwwvlkv9TDLt3RI8KmGaLGhaaO+4Kw8jESIM1HXCC+pdb/yAN/ur
/xi7Hw6bSxpXIX2tZItYQ20RQFtRjasaxzU0K9Lk801N4S4EpgrmZOmiBF7yNxHgT5HRp3jOg/8b
uwqHBtJW36PDOxefS7UloaFMCfYCYNZshEH4wjqP2QpPyEl8zCXRby1X/ffdPjXWc83StM9H/GZv
DHp3dYUTFhKljTCul5BtQV1gmHRwJ2KhlyB4tbw3IkdvQZ8GaIZ0KDdegn+FIMIA1ubv65W//4Ps
JqoB+QPyvkfumYYW1c2XRh2xoK4rXF6tB8QXmu2xxa/DWJN4j1tpb84lO5JKN1Fning8PzQInmJA
JaNe3CPzdYdoguBx6/xleRTUJP2l00+H5xdFOsPeaqd+gzyJkNufLyK7euMLzVRVFj48YgD3vHSo
wei0whxk9pbIqoLXFnAjQhhyMhq7rMbPfseu30OrrbdE+K57Nxktx6KNQ92dDCt5TDxFVfJgl/+g
3lRFE/SuN1kD7fvTHHFeoHZRfXNrNDvG+1gcFHs4ziHec2iq05lAxz0x71d5SsZsvCzliEL/cs03
MGOpES6/BGLiBmUl9rzeK063qKpLQCTUfGolOqd2kaUzG807A/SnD7Y0tcaGrSShcPfnMl95VL6k
FsRerTFddyDS/+3ouEbb78OaG2QAFdBzqabSBVF7KtpEdmWTliXaEVjOWqZLRPssZFwk4+hkwzBK
OcdFWTQ+vakXflCItp9bOneF3U6SeDzWQO1N6zku2gFdUaH5NaJ4EAEBhDIneXdtdmdjxunBZEA+
ixMloxugSyipesWC6pyuNvjoc1jDu1vkrEb4wQKeANJsUj4jx8peLJhB/LVQu5VxlqefOMoXWmW6
VvfSfrzH6y3fSm2Uks3v2RSMeuySnTFxymCcs/qcl+NKmhfF95LzjpCkmd2NUHlYspcWEwYbHwGo
xthDqD/riAmPMEYweOTsd4StFT+HJxyC30MPCqMFYQl4yWkqGdDCTFjQPK8mXiHqeEchrIhMZSxu
hhnQE36zTEHmOkZbqmNHcOTypAbz6paazBO/3TNASKHCo9ib431mdV3I7eXIPKrzv2TdxckvHKvm
LX7RCyajc8vtl2zlJfO46n4MzzOLLwNuJMGFhnt+ot5yMaDIlljpTgQRN3Y3PIui+jLCt1nuZfo1
obNWmk32/ntQTM0cglf6jqpDBFcRs+oHRVVqL4wx/CAQ+dc0aGpYydWC/TQgQkGUwz3T/XosQ0Fd
m+1XuimayKqRtPeHWVH7kCU3e86GkuZrdJv41YSJUTsxJohTWFH915jDCeuVkXrePzQzmX1g66l0
RLqJAOUmKEn97Oz+RPzwacMtLzU8S/bg20o+4dgIWN1Dbh+kOmNbazY7hcsXLKwr9FSE7ISsrz02
KCowXPiRI4jaujnOu+UkNRn4xWdKLo0+WCTgCS1WdlDmSfGeqImE1i7f+hRLkk1931gAjAkzXUhi
MS+p+9dqh8EooXq7bSjddOxmml5VeJbbcfRVaDY9YWodo09adZG5yJ+EOOkUZ4Jqpo5/lyfdRVyT
oD7UF2izoW9euA2z4pDQyDkiVyFCwgh83CkQq55i1/VCr7+jdW77hnecAA6g5hmf6CiDFgB9c1As
QXH35p0udQDIKfVRoypPhVeD4G0SJrXjAJmV7MK+EyEPEnJgnlhjfca740My+ynrBOzgc1jPHqjD
WkiDd0jxBM64NKYYhApnl6KBUymqopYlM67eMebJRhEFPvQtdHb47+jLl625Zenf8Hgxogklv8au
M0Q94JYRhp+zvw0UUoGSqDBNU6bfCO0cvlkIg36yw2wYXfbchx+382DPCqqn0MX3ZgBJsUJ+pF/F
cPZX2ReS8l6N0oK3j6jX6DWTA9eKxkZb8BDCft/yJfNgcYZEjtVoV6YQhtSa2IsRmy6X9OC5jd32
brsc7HPIzfsGI5asUUHYv562w9MqRGfTBzmCdvoymAC13cjDNsUIyxLK8nFIlmZcXhN6q+seM6Qi
nejvxRDPKwprC9T8dgy7Qadyt/gd1cui326sbvAfDVcoN8Ocp6LE1m0kVegIU2Qtxgly4C2H9Bys
ZYzhYgctAkfWYkZCkITdp6/jS3L3UzP5jqy3NND+5yZixNNe7LZzbVmuJ0s6ozQJnxJpJv0de6t5
Qd0BZ+sOSlwHK8fSTMAPisD4nLbKOuH4NjMxnYoy9IvRhBmi7I21nG2N12GD/I+ZgvWHtsffljQN
zoZpWRNPj6e0Bw54PL1WL+t6lEkHw1lBcWEgar0p3su8Q1ieCLs3P6SaY9eOkmWi1QerUBtmieHG
gIQrTFSnTdTLmBKfPnHILw8ndxCRyAQ5CVVwsWtCMwUZClIVBjGs+TQ8iM8DhbatXl/E5LFMGvUX
Ak4RuPzVdMPY4K4JDYki6yXcBazNETYxUuV+9ewbdhGLxpLG6+wEVQvn+tHXrmVD6W0p/e6ONEt9
5MdMAhPPmSsJCAXjF2VCC1+/55xdN4egVa+SwlkW75Lw+YZZ8AMSN6byfwrBE9T24vHKprd69wzp
1KgVpWdxzYUdqHxYkEq9y6L//h84yLf7IFfGnJ+VZJxHr4tcnVI9d8CR/6NcAcb2dG5ZXb05rlAx
1KXVopKlmLGUJTMMej4cXCSPE3RMmhW0EpqvmcbnbBV+BYFtrij5mGoqSFmVOjEDvNpww2uHoJIy
i4lEsoojR/ATlAfiyfJ3Ea/hibhbjX02CQahY+zjpk8v0kXoghNiMm0rFqaZasuBY418AWMXkT+r
mkz1Td6/saGmbaPkl9sfjEs958ft3QFSO09rZAmptrdo8BZca17iS0MrXvXQgl6jYlHeqISDbz7/
5CXWk6LAOVJFqBKsme+94wsaHJ0D9VYhvc4ryf9sayK8XAjMAapqaue2h63vAMONr2tNtJ8SGVsq
bj0Q1kEcftyg4gdofDapKkf/lOaEEoKQnHVYpKhiT+AzuO7Ic0XOS67nqWcXvdk+19AbwCwx9tGt
rSbZVFGXLcHdtzuxdJ6c+OpHQgY1O9rqtUo79duWQjEHp0J0M4D5wOnGytjrf3H1OUPNIioj39hD
UgZiFUoD2ZzsNV7/oUz+gcYX3z2TpTCHnzmNHmJBLKP/RJy8wcviZRHcUIuiFM3wNM6VQqYAVG9d
GEPojAkuGhcWnTGloQIMSegHuwm4zw/VqIqG+Uari6a5nZoJRZO7sp2t3pgH9Uw4TsSBahlJ2Uw9
AoGmd78h1dODbKOgAWfj3y/IVhnDtaHWOM9yDIDHmbXuewJYN2SNDD0yFDs9zzHybXwWfFTPYapy
7GviOfOUsNPcjX7aB5M59w4EVDqPtMA8PqwfHzfBv9X/zac6384l2cJf2Ff7h1YB+oYXTJReJBvP
4MJJDP2O9vfeheDwD7SzcSamKKeHvDv+KyPXwIBoTGh0xVrka5DgpZEszK2/Eq+GIhSJi3jcq99O
bZrg9sfMaPvgdD8Ndt1p71e1+YyXPSME1xNIIOPIZQskJ8n8cucxkbrDqzROFC/OdEi82JbrJE4b
WE7E3ubHPrVhLIBa2YD4Cxj2XhvaC2CT0ZHhOGjTvGpuhu/3lCTxQz35aqJDQmF1z05ac5KZgdnu
ehdwB067isnXnDHPwP7X0k4dc2aZI69cw4OnT8eiv91+DuGZcOMsNRvqmXL7kyuq4HU7PMvdJssa
HlcLIISXwfWmWCPnkqtYIwyrUrjlJ6qLJTBIPD9xkE27N4KKfRwt5T6s71lTMyWungzp9TbLa9VN
jNCC6/BDL9XI1Sey8yAilKFV+6/KzEx6UJWf3fotvR5ED/M1VAFuaCFtwQggiDl5rStPN/GzANhY
aq2RcIZhlv1sZJ/xqzSuob2E3NUKBTPiZfQvBHoKESJlyoiXPAAR5cN1dKjdlqFBLZAJ3PohR52M
2qDwp7DCl6l3z7dnmryCS7prlVzRi1SgAqDaJ5y9DtMnez8gsiuQLFmbTqjufDquX74INPUqFh2m
NCBdXob3GQD1tzfR3f5NUhF2hwQabEEsB5LanyJqkXLGZ7ts2TELKhoiilEV4TboH0ZZuuqFslrv
Nne9iFNTr+eJiNNIAnEjYHMieT1jYMMFSmcN831piHD/AVQ1T1TPIRijuoplB1FkNO/X0tjRiUgP
fOmyjaS1GsbPuARPI4ifAxQHNEmFaqJ351ylxpysxfC1IP/Cvmn2GKez5Nc6/9d2lVvm92yh2NMm
xHGsw5Ij1Whk1d38AoOdT7kCbTnkuEx2S8neNBr/Cvq7KsfhK3/fByoNXlkMd21GbkwkNBSpnOps
JAuMReRJjbqIuh2oS52D0k1rxHJzlhi0W2mIFqikDkOSSrPtdsE58Not+KGEwIVwcZbMKXLmjnPy
kJdSF86MQznduZbgyNW/wXJ5cvnMDt9v9fU/AJqAGObKXecLSLYB0pgvqz7KGNNJxkeedsvtBSa9
jymUzFbrEmFUsu976JUCGF6fTTb0XxIWKdjlUtu0wjpAGt7C88Pyx6HVcYRhmIIXHp1ZoAviRHAg
0zCBCImmQ7PysbxWXIfiVzfdsPfR8ZFZgo0mFDsP9DU7RqZOntqCdRZ4DOhcdUWsaO1+kHdEEqOX
aBiied6cFPXz5R4iAwS9YfT0OWamFSyrI3lkC0dmtNQ0pE/kUA0cMs3UvE+Q1tIB8KqBvDnU3+Kf
XmD8pvQtIsNKoy3uc/f1q3dV8pUaXCVGoefu9wfsY/iNG4sFyaPCXImSzDInWiKIchreOgaPvtKh
yLwbzwopw1X7yDfaO2fBr0RpuOR/jMwDWb7YH7SV/LJ+Cdb3n9F11AEileGcfWz+L/Qom+VQN9Pm
nQ9rcATQ+hJ8jW8AwoFPAm0spfy6ah8jtt6nOBai9BTqMvkzC91l2Zp0C5vOi3LDIkWwW5WEzqu9
oriblckWr5jLqnwedfnMWq6XVKVeSZu28P74oT/P7nQxZHQ25Fv+LvFQqB0V6eC6nGP0StKKZthK
VVQOZ7f3EWAvU1jmw2ZkyqgspA3KAwHMMmbbFSbAeGgfCd6cOcMsYx1njWZ0E3F4ZbgGf+i3ujJy
9H7PdHN8I0QaX/sNmQqUhMG/R97B7+whpd/HxnNyVxlDezAbKVZXliRP9RMzk/lIhmgNrqJ71L5t
eeQCf93u5mRX//WmiknFs/whz2qfvKzzuSHG623UKtl0F6Hxlc6HcXFeCp6lGCm7HCSEInroXKLB
WRXWypjCmGj9C4QQv325bHLfcQvU4Rhn/30HGZ57rd8DGipWXt98aEIw9CrImN/n467zwa0XS0Hs
ycxKtiQqoQQ9PU7/Yw9sU3n21R9VUPvv7idE9klqGK8Hng4e1VOzKH/tqODTLWKYoKsnVuyvmjlr
ytvQ21uvNcATW9JIT626B+qg9kR74PyThgz8kEiWnWSFn4RrTXahnegRwvPYHGAqf9sy4IAsL1GY
VnFT15TUqVG6RcuJsJWMIdHpgexuh0zYu/4ujooiy7gLB6Rqi3zcUe+w9x6ahOZimn8QXJHOQcUD
6PGrqSI9a5HagDrfjpAqHKVPPzv2yM+mOQyz7Os/l/0+o+bhDdDaaPFP9HkXodOvxYjH8engO1JB
PM/C11OO61pEyZBmWPMnJP6hv73N9PfTaguSTC6G8G5+z2/6qO/rlIFVVq/sNYILhD2KumG5znPw
aSonGpQnvmib9nsV+beecEcTxQl5yVaBA+JZLNCHb6k2NcNTZkDkicZ1wVWFSruYg6cU3y/7IKcc
eNQQPcAFSqSO9h2BmICw9+CDVOiJaWUnI+vbjG1w082rmBFeC3rjL39w34z5avZqPvGbHRNHkaOF
JS+Ne5ULB8uPMz56jQ5JjlRwWbcbJOYwBFv9xdgRFXTlhOISd8aozNA5Z+GRhsp8oBWQA+WktYvA
5smsDiELBdoqY/IXYWdINBvbo7qP8R1FrarBuqqpdSMRk8Z4iICpuXwjilyFEgGWqCfKBGPojwh5
r20ALEh0fw56QUCC5vAeEQ7RSslsoFf+K1Fonm2yw1nb38Ow9ZE50Vz4bqNytH2b/M8Fjq7VEJT6
MpRhU/Oj1Jk2f4BUtIIJcBNN03Hppfa+NEStUE9k9mpzA8ZBO/23IxGlt3ddOzzJFbdkL5cUy6ou
hB1PMvVEkGfSeq2gbrFboeeglH9cX0cViI0vdy+au4Lyp+i2j7bA8kz+ZaCbLwi+SVWIW540LBWG
H86h+FPFpSz/hMrms1CkSPouyB6A3S3/kHBpiyZvCgaztOlREZj0Y9+foAygsZ3It+wXOrm94ppK
1VP9/3/x6EGIr7e2ITZniobRoBJzcc18/WqleNdfjJrfh6XgmHzOINYB1wE+klwP8943u6zlByt9
Nb9pwsydryDO04gPGDvigTo/2mhJwUasruI9j3Lzc3a1y9oeC0RyzZZ3bNRMIH8nMsghkA7tNdWr
8kHz3G47SH5GMQaByWVLulvUyGdy79c2ubsIWePVqmk2R4lHEyavxwNXnhToi9WPRETx9GVuXq7C
oTIdEBQm9Brq2jcnXyhpDnaejgLBAte6ekPKit4SzfapBFxcyqX9dG04EhQFkg3GT/4JIvJP8A0b
LQbO2wyjxSqgjfoN0hKJ4YZbf9EMb/qTYsN8H2e9U/zhGHx6LvPyZDOG8Y5+Z+0TVsDCRMwqweOT
GkneNiMX8Nt99TtHG72E3OpejX/LZf3IHHJuh2dNi6vvME6Ljiuw5J2Fg7TgS28Y2VbwQ5/hO6lq
xy7FOAIWen50baNIyortQoAFPxJsRKE75oMJ6k6HSZ+7IKTcO4CJNMhy7pXKfwtNVpysal18pkAr
BzIX/IpJ0Ap42WcYHLhv8a078S6ufCwdxlqSyVPZsgCnfPyCmINJH1SMzB9LbClwXOo4+r1vxqnl
WzOx9L080wCtXc3ZnEaAO9yD0bl2DX2SNgXgdKyzZzG/KAyUPHP1BH2HPE6Vp/UHL8WSn7xGzHLN
Ly6mnu7xloGkijkT4KSfhpHINjh+vdToqb+6zbvfZWtC5HsNC1Ks7FzCKnmDDA6BfZt+ouG9d+U+
Hxek7GEJ81IabC06CUjdBbTGpJZZ2cf1AgmcWrUzk3E6fTvNrKVwheeRZsjSp5yjIMlDh2//TVMt
BjnNywpOyJ/x5+ch4VLuVm75w37PUz3+lqTdq/gSrbTqAGr2eGGmqphf3q3HopBjAI66A/CCDozn
acN0q/o/SEkc1iOyhgznCagpjR2a7/6VrxsJBYRilFN6Xj1W5BunPluKwIFn7QIAXhv7wfixv1Ql
a1h3JwOGWmluTExOu7+uYfSJnHn0gmzwiKgjgw/j0yLyS+msuUlHKuvrtbtNhBTf2q2T0QFFBAhG
RhsNTGfjk1nlWfluSWtF1m1XiUprs0KyrGadUPEgBayygDF5BNS4w/ucwB9cOeHvhm6TBsOxP94d
fVZ2RYuRBoxito6OYnp3XL5L4fAPAjx/hTQ5cRKYvHKa8LX/o44qItnsMxq7wckbQ6zEuKIir/nr
NwI+aYt93PaJewjq4QYxco+7pU0CxT8HquryRZ2b4wCiy2hzbLPDSFjpjr4+EBknjBJ6/w4wL/hE
bACbWIhhglpYWbvJnLGV3Bm6zxpgoFVkjBqEXdmDusXwaMTodl8Hy8ZT117O15YuppEYUoZepYfu
QOD4PC/RjCJ6DCL6vRD7InS2ZY73KR1kmmkF3i5kYTGrUXnT0TJ7K/Chyp1bKjTbTSW1ZaasBNE3
H6xq49d9ewHoCTtZ5ADL7qORTMm0HRgz5giC097J/U7Q6KBt0UfmktBcz+lN2N3nLToJ1JbNcDoU
6sKiJfE385Ok50veM5mUFCxiFL+H6KgJueovquC3pztFDaBLiu2F4xR/IPHn+4QmueM6C6+iBd0l
GjXMnICm59gyCWpN/OHD6977IKWq17Z8MAxj47YumDKu829M46wgN9I0VgrkHjagpI+D2ns6rOaH
qe0i24iswwJMw5sVWSknhVhoKogvUFoDsfuVAtfkQhJxso04SfCS/CC8Wkpa3siFbQvQ7pbesWPh
SQz8RziasyD+UjPhwuKQ1fNKx6JDsfkNFSnqQLNBfB3U2h+/lSPv1rl8UMQ4ubq461UrD+J903Z/
EOak47yqc9NMBpcW9gJxL6eJUYzB85+3hYvddCQV1etMDVpBrIWIHPGASZnMDEbkunOdILg6Dl4v
jPxf74mGhh9TINz0D3aTUpyfWTfeM6rcMsEWYxWN3Cim4XxMCWsavfZyHd5GVbY0ratkdHoALbfZ
C7hKop0Trhdr4hlVB5dI6hAsjDo7ABPddW7ZMTk4HV+R5szzMihNp93UmK/yXevluoY68j3zfgO+
468amJ0O/GnKL6w76dqMxR+rIjfYYoTjMyM7PSOKEDYtTTwJzAcobqzUI9sq6E4yYnSEnfb50Unl
TUnC3EhsPvupjp9e16aK8W+PeJalV7+4wR7bQs/utDEjlevetkUfULMGLizGTA4BIiqqlVuIgPtX
FYTlAWEwPwpRhNGOrmjiizEIcBB8BmFPTZp9GXq7fiMnJQeHq/3ij0SJgcU405fH0yMv39mahb3T
AjqY/Fc2MdqTqH/ZW5AnKkuOROkk5bo54H1cVj3LKyqEV915yVKStlnqMvN68tQM7UYyFTY2/aHZ
a1+gwgF3QHAbq2XV7+o35XyrsFxiS2lwFuPJIt0o0Hs6bcRajzWinI1sIkSEEr6cJDLw8Lcil5xg
3dlZ2vRSh4w4mYtRrizRTpl/p4N4fTRfr8l1TDO0FkW4kRcFxYSfYEJbpsDeyh5Wcjz4N1MLrJ79
4/K3H9xqfKGCs1PyihLTG2xcdl85QCUTf/IuVBPW10k/42cTh7eX6LraCoAv8o3Dpi7ZnnbVMMet
8QqCaiiSZf1wYb0yzJCc+1quOr4H9qnF8uV1+GFKMzPxuMuR3AQQvH5fFZafHelfxFzj2iZqFJg4
ihuwGD3tKQeI+omdzOJlaOP1WHIBNtyii+LNux0jIGqFO1eDW2vt9071QJOIZAwFU5x7aOGKa1HD
LKFT+me7KHHO4bQVv3dlXru3uDHadwHnEMv2rZ1pZdSzmz27LPnSg0xeYkWDVzuBtWxY851PJUsg
zsuI/xuGPus3lQU/w8OazhINbONNiPn51/4gM7qSnTLogLwPkPcfr9c5Clmm1xHKWzwcImGivVAD
LXCE/nvUF2ZzFMqNJN8e3sAQa1YwQL55r4kYhn+G0BvRAhQw/Q9qp4jJeSPQffvkxYrIfWduBlf2
m33Kw01Kr/8LtKIDTTKvaQz5akLIGibGn3QpvvLdjSTl5AxPgELpa8V+hnw2GGYb/XHDbGYXZntW
zUREtQMF7oMPhq9aCHtnzPBKk8zJtAYF3Zs1sdMITgKM/i6ddFgHqLgRKJI7QKSZVgXGubd3t1Xb
HUMxY44fVI/ta6kmCfolWELu2a1IJK/bt3Vbbp22TzLUQ1vwCZKpt2UYf41J72rjOLT+mfxXKqo2
UhjsikXj+f9nqdG6IcW8hOUPzJYtZznzlOMHEpHOXQJbNUpOO64zwTjpFcm1/yIf8uEGGZnd/FU0
oSkYcuxBR3MhaHs/X1OS69Mr20ZckCouGqQY3yC2U8CAS53r9ROJ3MVsAncAFOt9Z3NaFLU4KKBS
4p8XeCeo+fMd32gs36/eU34IQmAElCzqpe+oyvj/R6U/fy8qR31WsKzJj4CH8bkuoTmXmmcZQoBq
xJEOJJ7Ia+2hjEAJL2o+2RbFI/CtE/8wWkm9H+MTGVjvuGw6muiZ1GFYTwD31BN6PelCeAskDNDl
k+In2Ae08YeU0r+Hdk+PbszXhCdBCMc1/ok2FA5+t1tHynM7NrH9Ed5oBgYTs61nCDBBt9Oyfxk8
YCDdq5aa8TgU1ylD1wobK51Z4nGSbBD4X/SDSQUa0NBqpi9LeDbYfhv5NoV2j/yxYQ5dLP0ga8jK
TFDr94LhJXoonlZnjDB7hBHaV9FaVTy2oVb81deBaxePTFVJXZOQ/CcPNsWS1ihi
`pragma protect end_protected
