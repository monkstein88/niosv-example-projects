��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2i�>�|�"���K�W2��;#��Q#�;%�^��L��ǣ*��+ѷ�~ϵ[��{"��_3 ���No�NvHfH�E�D���;0�:5گ�鄅�T���σ��Sd��|ƴ��#��]I����&1�D܆�6�hi��1=b'�\d@����iW�^=�y}PM��~B���}5��Y��������8����5�N�i��y�V���f���V'�(2.J��ypw�]���w*\eH���lt���[L��s���ܳn�[�����q$�.\����Ux2a�.Vm�o�
��Hi�����t5^R���%[4��~lHT���ؙ�<n�	Ӛ:��H'����0�n�x��)�iϪ�xG1=���>�}��~6%�)��Z3�E6�-|�2��$Ұ��F(�!����Zjʘ�>uZ�&�����D�1��F��[���|=�d�G��C;�&��V�.��:��a�����7m�@$%[��-��\�P�i� �|?�X���3�:7Qj=�����`����L�}>��K�>��ބ�8o�/W^rs�͖����Vv�����sH俀��߆������8�w�p�_�ͬ�#)+���rg�)��}�Q"wLm �Va�*�R��R�Eӿ�	��^����������6r2��|���oY�0��$+�� ��2�(��[X�=\�=T�MC©81MÕ����U�`ji��h�M�&��zz�e�V����u�v������k0(.)��z�d��,�)�h>U�Y��f���)�5��h�"�8t��c�.Ў�&eQ�pJ�˴(rov��*�Ypd��X�@T��gP���ק����N*}8vRw�!��L��F�h�񨰜�WG�''d��?���E材� ��5͜z��냦��.��r����rk���KY��:��4o�?�_:,�ˤ