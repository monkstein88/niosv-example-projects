// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ucFmRTwBFwOq7qmfjbKszrTrjWXf6zPCG7FS/+b4Ss3lRE7Is+JWRYwMS4k4JxrcT2mYFa1PVoR3
PQiKgCYprS4sqceA0ouK38IEO3FAyD8NKneuJhIoIEWAp1jCOkiNHGGpMOO6/9/Ne2HaFcs4AIEF
5CRxm2/5KKcttpdxYYDm1CjMrV6NAM566dzSZfzFaIZjPUrnLGHY9iUxM4iuopENn1ZxaByX1zgG
HJuDlTjJKP9BFmK84x3ifY30yacWKk9C5nY7k2ffymWiAmypjpJDtwpXo9AAjTdPlFkzOPUWKO8t
FFg/rWAkN9Lil3JpfAjyadmrMccs/Z+CNeiRyg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 35808)
WimyiPq4IgriNWOR/yMMlQK5EisW1AOWXEesFXUK5RR+Cmwh+TczOEOedVmZCKj2QdjqqvZ7JNwg
DAE84Vfz0+rdMY/1hfYv6EoX0PinW2zEj1Y984lJEwaZYdQyRmCVkHwQM5nRokkr3rYhrb7s7hMw
FEQsQ50Qhiz9d5eLlRt6DDM0newTCA1hkPzvmKLG1BO/0bHx3CsrqHd8pdQh/aPLF47yF6K50DRe
XI+w5UYBpO4kDzbFF3aCAwHOk/Zr1FFOcSAyY0DSF63ldvwr9WCHHZ2GusBjrKE4w6t2jxC8faRX
JSAsB+5e5MhbcaNtJaQV8yRXvL067v11MvEZY/lmudssQKARKOshHtDr//IPOO11QWuzFPA4LJpc
/LT575eigv01e/ooFnXM7WShWugppjHfqjIZX74aRo+ZuYP88XKminBjdPJkDEk/Br7AhTmcz8N1
NGBZund7u6pl2QUvjdUDhgNlf8oDaPwcdlUJkzIwKwYHf+E/3SG/5pAAQjbxsSlZbWLN3SFxvb+w
JpGgdNo6qguZw3+VGyquuVYPk//ciezjmDRBBRi37BF8R7qmzjEL52Tu/5TqbyryrcJkcTjYXvdD
YbWTZqZhUYDikuOJ6XRDRIWGiS/hHaB/qVZ6GdQ5LG9vMMGvPql0xtXYOKRn2/u/KP23xcDzAB8V
6sDub3UV7zVz8prvr5JBgqfOW0eZ61+GpcSCg5v3z8bk1jZqwjF7p1O2gMOdmsF05PyRJribxrIy
vkWzkivFzIt+CXft+PwNOc3UxrOt+Ce9Pg2CVLmleFQ3N/ONAvLT70ye4Qz/BbYsUmXakqWpfSvN
JQjaa34XIyKX4vuA/1Cj75WiGH7QOgcEPvxzZWJ8SvwfsuSWXjLg0Bk8IuF8ruSew04Ha64wZ/S/
Ggxp5p6oyVcgdqT8pS3cm17k8FLd+cn0qarUEqSbSz01+0F1ZmvNmdCDYpbHk1YA52+C2nzq5EMw
gsKcff1U5WjEGO5AYZGWmQ93RoOOyhR7gDfc5z52q2gcOzPDNWIegaVlgZKJKwIYxk67y0eKeJxI
Xg5YlH/UAe2FLOR6laqBwH1f+gWxLRWkwPgKUHSp3V5UXfhaHhqD4SfS4zXd4RhyGkXEmLqdntMP
GOQ0kBEA2ApQ8jT8bQgMWNkRkOv0UQ1TwQSiR1lk3IrLrhiWPO/MtioM05UFj8+xbHyUbwCXiinu
pF/jUmzc5nuwEtWGPrwCIWx+UcYvZ26ql4rMlDG5Vilillw02prel5xiec9r79GlH7RPxoD9kgXE
NNN+H/79ONmM6fH592tFOiMKZBnQKUtsQ67T8MMaOwEFJZYVr41HQ7LqWiBOgQEi3SUEUtb+6vX6
kpyh9PDufVAhTqa5K9qH7g75tB56gvvvABewzU3owsRrpWw26hISH8jUnghhayQfOQNlzPCfD6hq
IeWTb+Qlk6DCta3lio5GjTVIYFKQC2cMQbmNdQbwvXUTInsDy36CcfqcvecSN5wJXAO6u6Zr0Aiy
tIYGKz7bXrjQhFKeUle7sMf4rnVBff6d6mwfXrtVExQGCsoLIHXv+3Tp0RA7DTcQMpnDbhkR3CRl
OWGqLkT2Io5GJgfB06CNzSW0PYk9nWDSQk8YZ7tMvxlxJPaWFYjjhifXy/2SSmU6iQLrarXvJyJR
rjZB8NcyRR9ETnIV7QXwvL9M1Q59U9/nLyzG/0n/jWebjtmreQoPaD8/RnKt480rcAGm3RTVAk+7
vsVZg7VfLI4blU6QL/2Rwl1pgGodAXCPFo90BVH7WSIbo8bo+t6W6mxDMLDv3AgPLHs7Kq3QpNo9
BmwIWzyGz82JYcurXdEJURMywZz5/pWXDIgcmauIWeime8S87EE4fd8Ny66xP4Bof6qqXtt8AhTy
7Jdjpsz2MXgNeRPEANFE7zIsqR2/xrNZh405hZrlxx3kWYd1SMa4VbsEgf5yTbAo/qBR3ENDYOwF
oU9w/vA9D0mH4sUtVOStmFI2G43AQbLiu28tN6P/HAmO8cMm+1nYBJ92iAdm7OPVHdgpGjITitkp
+9axf1VDXvVtc8IhBpd4Bjg5jIHzBnPV1CKXivgsVSQtMpGTijA5POgMGxL4xD34tCFcCaYB++KH
631QqqCPQhVcA5SU8rQRPPjMJ+Jt/P2a0W5v8RdEumI+nk6feH4U9rqvTcJapF60ycqePFS235Yt
wV2N3wFDHCt+QuGREUOxugdcfEjfa7ynkUsjkkZtNGELuHb8wfNvr4+/RsOQbo3pgQZJnxhq+8sY
z+kemQDCpb7mgVUZ47+iMzFSIb6hHR4akwXQ2SCJghChYWB3hLBUc1tTv9V4Rqo9snNGQupScbJo
Vgu79tvOdVtLDQPC8ZyVmxrLEdmUjYMhSXXgLDdWUR9ZBooA7+yanvczeQnNjaDvwwnn7onLgvbt
s34wPKT3YqqQvSkU6k0VvO7KczYEgu8je9qeALZW1tslBFYPIemimjpe82oaVHXi+tX0XQnuwzdD
sKXHe8ZS2js9Qdo1QxetZSD9MfkNJlHHaAB21OlhpDGZ6xwfoL50HYrtM1T+Sy44HT0nGrNX3wp5
WUaxW8uCd2hIkq7P4adOWKDqKgqRlaUfoWyZ+DGAMRtZklXgUvkvxpBy3/gbgsOzPc7ibGhRrJNy
uvOoJG6D7py9hbz/0oYazSgXnUNylcTs7C2CjXSyPrE4JbksrUfwB2z8q2b3e9UuinNGNJbaXCyA
569pCnM+KppTVUXUuQJEPdmAN1BbzwnoDR4ft88sBf1E/LenG3V9NJZz4/2ZydwtB5dwyO9xZ+Jf
HWc84kFifjtnH5eQlhtQmdKuR90aTXnMYxcxRBZh3SFlP5168Vsdo8N4tIjY7QLOUxXgOi3zgQm9
rnM8i6est4OcHg7kG/A4Dm59GrqLn0R8FQadh7EAHVIDFF0dWUx4y+8xblGtGP0yrx8T1ZfjdcKg
K+GAn/burDVR9xbmX2MhNFkpeUi86Tg8zOD52nsX2ISuC7U4bp2vAQ5o9z1Agmqk2DrhLtX/tqgD
0rWB1SP+E9luBvPyg3QtE3JiuBSNHCLZMpjFlJJe8JBHdV0OOxP1eST6S/+kmupuDys9p1SdhnB/
0k1pclyUW4jesN7HwNxB9M3LGqIJMnUGv5hfacGahaoxD5v7Un7AzQTguGy4fEcmWFEO19KvrlHM
YxgdGQJ+LXOo8cT9DfPEGf+I7g2n2DQkSdhseaDaWmVDlm2wKPQr07z80KmssFx0ZL03rp0wBHvA
C6wOMzEGe1SCKtrGXZTb9YsTsobRf8X6J5IOtbgi1QKf7E5CPQAvBByBZxqwb73XJmWZt+q85rnl
HBRPAV89nhbO38O8PtgalrPtBGNfmwO7pdwEP7WxadVA/9nlLotBGyEUJjiaRl90CNYXeG5H29PC
PwLC7jOOp2pJ2NEgDP+VCdCXBA7vcPtqDoFwk0iFKKnN4W5qUR21E9fvw5TnyA6SAttzjGUCwgaK
/HlicdPoHzN8BmddySGUO0rmUygE/tXT+db+/OjkcSyWehLQ3Zhx1JuP1y67BQNKhKT543g8fkLI
k0Be90sCywL2W2jigY6HvUDlcuiyvKndxPZBjUAIhPcMg3mgQA52QrmHz683EYsbRa8x6Pr8FS/C
IYUDR64SzeeHckzhXiRUmay+I+wVXXZNDrWPoWOU0KRRaXVqLk+Dd70LvHxs47zkznEpBmTluZVt
ItbvtJI6iAEH9BeSg2NHs3+wFYuLcjxbyg79nAqUJNuE76Zp01u3k24T+fLZa/yL//fcV4ePsPCA
ZW8VVUr+m48RQdnzueJEL4pVHFwNnpLkSHJPr4THCtpvWFYmlIS1T7/CIA8net+3PwnlodOOZqP2
GZVczJqOqHJvghffZQoimXp8VJA8Bv5XBpYqOayhDmmAypdjWXFHAMgwaOieRV7otOfYFOSQIjmI
BvF5KuhYiy8lexH/mXrXquFX3Zt2QFSflFX6Phmc3Kactm2Nx8SNm7WypJygmNDQLF/vJw0AOPN+
kWZlcXnNNCPimxsgkFN94SA46kcGW2TEQl9bKRv4k7ekpBo7MO9qc1uP6SHt4rq4vJvb9y0qjkFT
e/xHvwZ2eE+T4TDz/nhCRsJXuWPVJc1Pw8O+y/jQFmBhDhbYxWUUjZ2t7ah8bJ5WpoWlIHHqDijd
LvBUHSGANhQD5RhT/JWw2UQvTJa8YtmLjLmlV2f1oFJZPRvdUQh/Q2acD9FyaSeKZDBF03efBp+i
QdL4F2pm16cEbIMUxKi3hAckjUdAi4XsfBDiOzXOqt9IFb7oxJ12peO5Xgi3CXqTBrKLLZ8CKS16
zr2e5ZZFOib+dLhpy6IvOJ8jK4lJy+vSZj4/EUdryCE94asrIXOXMU7K15zTCW4iAelTrdVdsOC7
5NiAVVAcmOttRSpkgB0kKTj3NIK2HsPAdpAPCdUE5+BMmW49ofdQ/eKvNlAvwNEpRyL6udasH3PM
Oyw0vQlZgA5+7oYt0AK/TjL1sJ0BAK3Lx9ZEkZXkmgsxD4mKcbdcfionoottodC4fLzjvMygiIh7
FPdY0guEAXxklrvb/iggb3ol/J0XX18A1o+pZMn78zvDkECkAxmjVRjYTIlIdL+Pu6iF8um5WEns
dVsCv6/u0vEP/3WdnbysP7dwf+AcHj+jgSabtU51fRrZMAqULpnJf0gQzT1jHF1VnoYj5nyNnIXO
3nWkRAhdi4zCck40/4DmIOJuzHojT4balKySQS0yIsYwI4VzzXv6kjDjd/3qVA2wHm86K/1k8kTP
pDHJRs0iSl7m4o+QWm0H5zh+Nh8T8SEVAGRmB0cxIaEIAKrbAgzaHjv75UFD2GOzA8SgixI/QjJX
KleSOhPLykBxni9pERGA3dsMWIqxqidj42zImo+0yc8m65jEmepCMsyHMCm0E0UEjhzpc8shHsGh
WeBnXJ+guNRYWxmPnO7SIfXv/QKfduBBFk09pwqTHl3VnuUoslbiMD2DHnucP1f1gK423LDbL2yE
VoOAk7NVPwFxurfqh7jjsXGSw+x8Zj5QJKDwR5sYl5m1WaTafma6MQV+iLJV8hUphDFK+Lk26PKG
Rye70Q+/XY9dc90up2z/YQ8Y/wmGDohiJuyB3EP19kkx9tI+XxFpHRLA/EFUqMgtK3IW9Fl3eJi8
KmwXsYiAqgWzZ2f0ZjIo5ctxtTLM45Sci8vH45qbAwNEQ7h7up4URPpEzRn61Q2C/qi64XHCl8wc
0v1ejmqeNwMyHnbg8+Hba/hrf+8PNkv6a4Q6HBYlXnytms/EJMXgvJw+u3kFnOoCAYuwlS4O+s28
FArPKreTPDhUmucvUinXVd1GSWQjgZ78eCd/s49gi2i2Zai4Jy+qHmK0EAnJ19bwSXEvL4R9T/EV
jIw8IVu+rS1aAKq9/r4Q7x1AOpZLkRzTDDv6g7GIlLtx9kjTsD4mBqh1DPaT9LBBEW3J3G/+wcNs
pf0fECEa8Vm55t5DhNT/kuGxakPLLhdVQktDubcI8cO4WqLCKn7F60dAMl/OcROtBxKN+43MPYWk
k1t5hm/NUV0zwEI88zLa9vwRJXat0Md2X+mm0NOhA3nudiCMwAEzBpAxldlJM38fVvf41O3nHLiR
DxzLa9JLypAgw8QdYEGMpeS0GhtkV9UXD9+VzjXMmFhC6fAk6SosaLJmCdAdG1RDg92GmqR9Jxq6
Piil0QWEWv8BmNKC8Msi8osGkD/0ewQUlQGkZbKhpCm8H8s2QI9demym7VIDY1QlI7PKe6jWQhpY
ztYKGLv75W8x9sDoPTTfsoa/Tz9AJMhiRaT78Zxm4HtXNAufLQhohycaPe0OrpbQwyA07AfplBOv
spnHVZemsDgaJvm9v55oCUJVIm/53dIuktNPSiqwkl4U40FWaKq2DuwMBMX3MJ8iYmru0rAmz/sC
1lQnVWizOGhY0DqkwcntsEiU5fVqN6KTVu1BhbMU+OqP8XrXDrWHWl1JXafWir9VWEF/Ivk8zDY5
gQcz7Ze6lMGokDPgAnadKGzT6gWjlTNDc5NoBKsNym3QBe6STGv8+8KjvZJ3Ns/FyNQoNSqlOH7U
xcPZ2C0ySaemiIs5piAVxdnWFAelCioaGkAypwIt55MLv+AaXhDLfwZl6jL/LTV9xqwfkVaNwak4
pXYSkhPdzDD6FVvsIubzb1ziYWx79j2M/rt8Q6xaEsz5ALj+AdHa8IMaxaMkkS+e0Xf5+NhpRVoT
ZPoFjTsS57ZNWPhyRp0A4nJvRkyOrVY+XtgtIeZHdKhfB7lbSWw73CH9//7UUFUulIYKlMH0ey37
KuYj8YgxnL0ayMS85bzphPZfa9jAa/feai6SCQLKbYjI/8v3NVCUL80KL53+lvOGztebC5zvqXvX
WQ2gtSVw2ycwzYLaK6iBNoAm1/OSAr4s7H5vlnI8UHt54Iz7pO1euN6KzqGZQRdHEUbUNbzxG+bM
rFfMJHmhlvF4QIzMILOTo5c1Wlbl1rCtXWZc1ngHESZ3eglAKt4iVWjRnoOwAPwkNLMzNGaM00li
T6QJqnI3JfbUwVrNrMEM3ArFZio46NImGu9WS+morFp2K+cSml+joUwtWvzKDVq9gSvgUHNLmPzm
2pko0cRH8hJ9Dv+EUdubHa6aaKU0nQa+1u7cYxS9WuZKEyhCqC/Yk7vsBPj9QEscwoQxxXR6biCl
2rKdvlkhSlvAWP4JImVSX3vwD1I/Vf+YJTRiXtcd0owkhi+1sWAl7yM0CxUxrhlEUIKYnaspx2pG
CHwfU1Wekn6MZKKV0KhaIWz9MPWF7zUc9X0qC2fbq/8F8HFV7H4rK4S5ZTFMARPhzqkBWlWCgTXY
eYUOBoVBLmO2Dk7RHWcSdfyVLvoUTZy4HaffKREKh/NecE/gIClvj8NSiQGp6MOPFhhL1nR0nUpp
orPE3rH7Vyh16HToCJfns2lgwDitIgUwPg9nz6ye3/YJzGGtjpqr8EuvmkxMpSDxUgP9++oGPx2Y
qKEWLGQUxuSovh4bM9sogKWZMg4tqXCRgXYWlawB+YlNBIWcnToRnoWDQpQPR2s38hPSXUGisMDL
0ukUXVntFNN3+gU2Z13tYnLr7v1vnTWSB6cSxl01WEh7Hiru054MAxcmFId/2lYaX4ye25neIoCN
Daz8cNw/6E/vIB9IeAdwzBmylfOId16QQg1C5JIZHnf2nlegXiYv5gORzec4OxLAMuNTE6dHUgU0
0Yz/LA2Mcue70r5H/mdmPyjE1t/qKvAtuyD4ENKmAgHMEKqq04jjYLe2rusqt1z2EXD1eQEYaDeg
H6eSbZ/sc8o4DdZMq+2c2s5DUrY6hMs8cw79oowABpMfn9JbffflebtdnXH4stK/fcw0q+wKAISH
po/HxFch6nSFTeL2uECvgFaKJvsRqxTOXIzvpCFW6xeQdfC8281F67QxWioTu3ePclIYSOEVxBJX
28HSJVqtp7JyYsVQ7XOk8gKoFRgGJaYJjKrHu3Gk5LmbOh88uocFFLFzGFcd3aNNJMyxns5hJqjM
XgvgT0Y/PSLy1Tqxw26mOs9MlWh/jdHDFDFC8InVRtYkW0j+YyJHOcjzHU65B+V5XdkFxc9r9OwZ
X38iRtDT+6eIKsSvgJztNRl2sEMHeEGzoVPMA67R9ivVvCEXEoUi+iF4Ckv/94UTUlaUTd2kwshL
Fj7z3/wbebQjdR+LmMFOvsZJwKY+qVp8PJdFQPL/j/4ZRqVYNhNMLNDOTGIFP9StpHn8xJuWT2Jx
we8O7WG0o6TjeM+4dRCcgqBE8edlb6VOduVAtF11HWK17v2oU0/RRaH8qr6NHmZCoBNtRc6/zt55
JHbo621qO4+3YGtTJADAnOvRDOAp2V/usdi07bSsbuBG/zpYLRBUuKRIMWV0D5IsbXwT4th9FChq
ZEA7PTYGNaRD6B6iWfABrzlBybq8zMm42DBV0qcELBMnZeP+/44VpHAtX4ZpjtVMOvpVZtlQP8ew
KV+E+OVQfWEB3BksJKAscF+FlK45egPWuNawM8ygjT5yRFxTWRJjWRafyVPwMTVH8lZmrE5xZHqY
d9AHVHLl0OFBgNk0hijcPwZuBMcK0oFggcHSUk9PEmtIsOg6gqiEPeraguPaCidvKNCHitd1arIf
2qT3u+y2Obvtgo+0Q6v1VsD0sI1P9hiWGBLtdNUZrBPwwrsRjduMvBh4lNY7yJTNX845Ntu8YUxj
8O1EyC6itNimL60I5i7tBYmfIHUCmiuEhoZQJTBWo7+GPPpyGuncyRcsOqrZo9un3wS9PJXQvl+f
BsOYbTG07AQNnSmR9otflbUvIPbSkaIcmw4MhHY5cR/bDiSjeBWJtd7FxeZ3zVgLVNpfVNy/rEaO
rxjMvczR6J+CNrzefCLsTeV/e1xtDdBj6LyVC3/lXZmm55Jk/l14Kn9wPQYHIdEs7Ou8s5RLHSTX
bTRLeFBdb31m/mzuXpbbimkq4ycb37EkiudFfMgQsLdKgiN0e6Ul/BnPB+RBn7N1n5B2640DLosO
0QNpSKI5CD0mA+QhECWNcTi7Yu3HVoIer4LvyMvRTedetZyL87yA/BSVKWG/8wAkYibENRMiAYzK
A4z49ufRByC0DVtPXUzH/NFtVC2PgGv6wL7iPwaXWfeMtzhdZYZpPmts4CbqUa1IQ7ArUMSuBoJo
N3wxrU28sAquCLjmWHDryfJwgD3Zpdou5Dm3u7jCZIR5VvKJazuyN3m05zBg7VtxTUUPvAYIYuwa
F7P40rcVHTgaz5ltb+El+qgPKSv+BM2pINeZM/dsr+fmT7pmUbWpu+nQ9BhBGAbg/SX/CV/Sq/9N
YMCXJ9IiFKCL5MIhlHLGLztX9wWDdiWSI8xDjMOVgWRg4OGUIJXL9ApWBi820e1HnFE8UGjiKiJd
81KZ71SYOGENr+YytQhiALxoRVb0apA+FQXXFVnN7GFl7vjNtKlCi6yFYY413BOWwgGXw6xv3Vxp
ZW2Pc4TlJ6eb+eJ2ZX24YZGvUJ+Df2KubIjjvhsTIIbWKOW9tfEiKY9PnWFw4lo197orLvHU8XKy
z/sAoHFMkHKLa2lzlA0NYE3D52dCDcaB/dq67LDKRwBL6D5ChYHZsqmNSP5l68Oyz6PZ7i1Dn76n
Tra0rmpAYA4Op1JPJCwE/snU7XPe7Pdaa1VIthd26jIP4mvqHlgbtbwDpVvaoctgwOu+8PmwGj59
qGycJRShAX5K3Q4rU8epWuIOs0JaFfd1Jyp+CkTQ+uU/pm/QkAXLm8RPJbS1I8nsT9aQ909xtB7p
ssVfIQNXqOOmLetvSmhMK7VaMd5614FRl8m0UUNvQ8LJQ1vhLdJjP9737XFBMYZLJbewAwIpfMvR
Hm7ovOjrOucx8d4lTDGTuBka8HFzxOD4AqFBQqj4hXjaHNwZ3t7/rcKvICsybNRaTWyeTj6+ZXUu
1CW0Y8+dPqrptW379cULQb36WlOjSFLz82OjGFMuvM2Bn3DZGMRzgdbyI8UJJOAh3pIK3Q5m00ep
7YvqYLOpf14wVzVxlpenmwmTwtkpNMmkEdM6i7KxlR5lW0pvztPh3EZU2OnJMKzWVwM5RQScSCrX
uql99iIe8NWUNIN81HXA5DbKAyn1IeIXvIQ7cj6BjiTS7XzmvVdcwaZu4Cjwl/FbdmkJSED2CsVR
S333FVqPXm/n4Di5BW4Pns9cLM645Z6bzH+orRfRw0gsr4cfY/UzwsZ3/XEmjPcSVIxgpP6GTPR6
m6fwVCzPpix+sgMVy5nYjKe+E3K9uyXePKZBk4SondhU+3VxMlqA4wmoKYcedDy5txHG/2aQ/fpg
1qX6kkOlXiX6nll26vJ4IxLN6dyu8av+g1nkQOtjiukUzWE8ZdPBcR1bBjPj14TnOzoAHulFfx+U
u2el/F/41SOkSUEc5XvPFD46mTT4xQQq8pWQwDTQQPHlctYWM+aAHOAxtDvUkOV+ygN9XCv1zB20
/ecLoF1ITOFuGs6tGIT3qZnyH3dK0iAjVsdjhfzCjOdRdvmERVQPbcdJl3brbk3Icf0xb8jCfVPd
QJg4EJBj5YRQNj4SyX96+mtehLSyLwSGaxvnOTS9GiAarBzUcjN0HxVprbYNmH3gxzNXjUohbKue
dm93ZwNo8jtWzcmEgEuU05SAzy6lgp4sVesGFJPwRiyMpZXuploxbfAFeww8NFBtJ3pETwDSh+u1
oF4elCwCLYTjV+OxkEz/mEfV8A3+AvIPy33jTQwNoNKH31TPLVWKzgGVzgFsQc90uEsMMUB/ReO+
wykTlsMfDuB9gMws28IuqZAoEqwxYjMMoIxWonuDCgubhTqvcJXnqalT+9DZmJcgNribk8/ZyUUr
qHS6YwQYBBmf0O0mSzPOU6+mWzxW+vdawXPvWusCumj4IkLLKL2j3anBo6IUNVy6muIA1tmyBH3K
alB5K4jnIRk+W9jxXufSbq6vQNuLDQ2B9oZaNwIXzNTR8f6AK9oNTKVAJBj9r936skuP12+GiqX4
BY+bL4R6OrHlN2QRaUfTnDQPprqei5S44ys3ircFO3s+9NNJHrSDy/QTsbTaRvhD7gBf/eyKmBiK
+f1v2lVQCXheNjBW4MEfQZ86aiB+nMWWkE24iEj70AIAyAEg7KdoduEVY95DeH1USJJpWKr9Ydyp
jFoTQIQe2kFOiOZWwCYwmctUQ38LiAtL178FuaU2LKh2tgVi738HcB56fmrf+boEmA5RpypNCnCr
9v5XC6t9P8fXwsRINpNqB/Dc/vFIt0oSIM1srN/2o1y04yUdQ4jA+WtF2GLfMqdNpmt4LJofiZDH
ynRPWid4Njt2uOGmOwx+/OUN7c+QQbtxcLkJPMIlyC0rhLYvjA2YSoqxLIjQ9Uo3iKDsQZ0pN/pJ
bSXokJYtR3BwN2CEy10BB4QzW4atU5Cz5Y0RGnSNYxsJ9d8A5icQrTDJF5Mai3HIS/+pAMeGtf4Y
YTJKLTM1Gju3XtM/onOWe5gT7cl9GSK0xt7SKZ51GCWtA7oYswLOd2fyAfYeJB9WH0Cmn6qFqRf5
mwAbGv+71XZg5dkZNtVKwfTvulGhAEqkIurQ1EQcpThMJ45kUBFOhvnwaBRy3mDQ/GC5SALrzPay
tjssLkjO8jZ3e/ZJ6KIyYiylgFNA5pIG7NS8UqH23dl29OFDovyrolkXIhdLX/OYUqMCItId4UL1
t06tN+R73gsbdH76UbQibaE2PBBsp83QSi5Kqu6kMrldIlADVBRTI5mZJQGrZNWEjtfl7sJ3yY6k
cRp7qex/2XsJDDqJDm0O5AtGjTaDi5djvYyppChYiPpCCkj6oPUAiqCKWfJjcWRTWYgl00KPD5he
0y+wKCl4LOOfgXRutoivSodYLQORyXgl2z0AccI2bYf84FMXOvBK5SR0MrL2+oxnvY4KtibfdfkV
0Bohs2p9yhELe1RFUZ4Z95yw350p5dhoaTazQl0kuqPZZHusTSJMCG2R2e2MOJX03ITrkg3vIFwe
DD84KyOoXxtJ18ZkFSxXF/rSkeIcIz2bEo3Di+gXNZuDd4NA9FEzlvLyGHfCafpJN1V7QcP4r7q3
94qBwc1K+WlUNjoFV6NsA6d+ub3pLBMbjo8klY8xhMIkMfbGpnyrg/IoCJGQF7ZbWl7E5Tebccmm
g3M9W3/59zVYZG1O9wPRRLKhuKcSTAnd2QXBzUQ972iUZV1lbKzD9J1JS0jRpWy/MtElU0S/uhbJ
UHiyIQIjYjqAQQt6Ab/5KAR4hRfRITF6+s0lLb3vQL6q+D1DcJjgVcAT1CaqqvQBp1iKRjElycvE
i8t0I1gZpS62vaAM1n4F4aAptzRf4zdv3OF6V73LvveqimQmN+UrinWRjqRY4afnL1COOikf4kMU
9cFRdtRFB3mHbfU/BM4VwL2nOvAG1urHsv3hyriJ53fpnzr2zs0mnskBfzKhZAbvzGtZrfABryJT
f/UKT3rOtmOdovDk5SorGG2GDG54+owAMpJSUiUHMwZKzbvhj52q6Ayim3SM+e1uVH05Ls9BXt1t
oHDWZY074AroISNW7BbdOIL7fSzc5sC+pMgqaVhSKEwBr2Qr8hMBN+ps22zlHUiEMHVbdGQR5HBt
B3tBJ9J6rOXnm7/AIu7pozNs6v46D1UBiFsXpTngTf3Dh3lrea6vF2Cvggc//IKZQ+SfZqQ1h39W
M62ZS+PCwNmxb7HpIwCK2ClY06qOoGAooVPU5nmIx308N1fB86o/mQqb+8Fc/0Z10yDOubOChFR0
3h5tLLQ3rtjcx7xMxin9wJGAFdPDAV2Q2dAkgk+/TewwHU0vjEUUrryA0tdZmcpt8ZfO91OsshZS
cfCrNMOgJQDBpFEXILCwtMCPruABZFj329vDam4iCo0KQcSI4PkYJyDZ9KW8NAXd2ULWd+A/gxNf
DV2suQKjeEpsV0hgMenoEfRE1oAyb05vvGPophPR6Z2N5CgqVZyWEhQm28Y0TXZNwufGYDhcxCT5
cTP4edAjF2VLy5S74QK8a3GDy6Q6LGDAZn1LdEV2li3klM4qUmrvLCkpXqb7S34N530a0mOWMHdf
kej/emSEDX9IruYaxuYRtBauTnzmR2VUVbzsmFQOSEvNa0KyWTfUj5mxQuxNjmPDpecyqGKDttJB
WbDqfPfCdn216vlC44dYIeHhSwoyJHSU4RHO8xgJR2Wi4+6TwdCOkZIM5LNeL0IzoTkiYtm9DT1A
Z8h2HkfPcEWmTM+nUGQ1bptmsGtYpPryfewJ01zNWUIiCoExhnc26dkZl54nErHNV11g1CqQkUje
YMDCqTUMnkoP2231fO9kqzp3CLiZhPLhiXncKJyffDdhpThUMG0/DjNSPXMMDKp+klZOYnu+pH+1
UvkO1BS9O/DRfsCYOfT6Sw5tIJ4MZXcKUNZutGHt3tPiLTkJ2YxPjOuefjJBM8SoUFAMjsMPnpFm
pLNjWCKjWf+V+Yj7bqkXQ36ThStL36mTZb3i4o1P7RTbcjBHAuZv94CiTraQy0xo7BplrNgVEZkv
A/+kuD+pUCO+nssA4kcjJK11VfSf1/0eICPPB0WoaX/+x2klGlgvFU5hEwJZ3qJCbUVvFuAcNUgL
NMpA2Xq8ZL7WIcffa/wLIe+6mTsdL6nY96UsmKAB1ZwTtxlGc3JM0E6vNscnTFKRYhEAYNwgYrH7
cV6Z+ExA18D9M/T7nbAA78UadJiKwnboCdTHtaaJKXJo3hY8jYpQcOECrBDsSZ+W1lifjhKy58hN
DhjveRPB5dGHuTZ0S3igTfexvVZr45twNHixJeAjdpGmAakA48iHwFa4XjTFOZWZOjLoCxbMry5t
5Sd9NPPvFdHnrnc8Li5S9giqqNo/4TycxD6A7TnldY8uTCpQkaiMWzz4k68IKHKn+DKQ77jVxtYr
1xQW9gGAYD9SgEyLjZHuiiqW7gtQYzSW18UcJPxHPord2TiICqVILUf57uIGamNkl+Hp0mr/Jpow
3KQ3VNs6WjvvnZuDbeQ6nGgwuBJgm5Mc8T7o8RaMIwVpcGxoW8vNg8A2Q2Izkx/tY4BPST7dAD37
JUvZ59kLDOqgnvH7i5HuMCN5CR0wzadkqte75Ic5aM9Ukat9DZUzg202OfCsyfDWhhhdiXDtof6g
4I/0Lb63Vja8U/XDrFGD1+hskqVaT8WwsWE7aIZ/qzXe1P7BepLe2nvbclY8Mrgli/Ds5SErsLcA
27XNekco3GksjlchP+D55BCWjHLboFGnkwzzX4rV5iZLG3l6Y37dBusLvn4hr/dMFqO6/2E7dluu
5MFR386RfJtX5zo0r7V+PaPWppZd/g4dweJOFcrXwn5Dn/Alju0J9DqC9orQAyjkRb3a5WD+1y5i
TMRNmLVbnxKVVrNMg6yvwGRmM5C/FZJqkCNlS+aYl4gRbcMNk5xS3bWwrn8oj6JM94CaMffve4Ck
T82sBvLGcce/TQqLdoC4WjJ7Edrmqv686KfdJB+xSOYr9s4+dLgOv9lpoNAFN3JlcrTnI8vN6QFo
V2fO0T1aOhnuyqOiQI0BoX7RQHWw9pb2vT9Lj3Ze/UG51lqKf6sUldbf2MJtMjDij0Um454mNwzJ
czEomJmSzbd79hIsHrulXvdw6Y4aj+hCkjn/5AIFEJTJS/0Fu1pimFWLJa9bsCJxzhq7WPPLknDf
K0iXBHvgM/aM+utCctBgbVGxgl2g0hh/mK1Cj+29dggKf36+eGRe1Nv9kBmwK8gtCSAZfCtxu+QG
hVijCqilDRCz+c5CFjJfRGsdwd72Ro79ljSXqwvAlt2iwXsk3Bcl6PN26va1bqgCRTSp2JwG0QYX
vpL7uubkxiZfGIjPwmQzIIOLnW81McFfJ2Zuh52bNCaH1wjSaCJJ7rWxoXGfm9i3mPnodM6qmE7E
9cNNFsP/1Xug1ECAJuV4a8W0Ia929WuLmPiDOQVky9yXzUMBKxZLKL9uD0NTd0qWKUpdWs4WVoM7
JjizvNy2W09aKaRPUALczMqV5Mwb5ZfuYcbgd99nH8QsLX2gQWPZXWQkp+VPcPaciW4adFCBx1vk
afhzYS2ClWhcbHN4lFrnlhERYVMIAD3gRScQy55qJ5vjKEwhT11jbD3TjurftHi5BZ/TBRgyEGfK
XV3E44OSPLJM30v2ZALkJmMfGkn4QyGbxjlWPo9LwlmBHFmrvsiyt0IUcX1s/yAvapLtdKTqiFrt
0TVg5YrqGspa12l7fIAWH7DO0ZFhJF5uao/9HOtxkNqrmE4Xyfd9bNoJDnd+Zm1OTQ/D/aOvzMpP
uUs4pWIM4KjB03PxDzS+jWXu4YpHfWV1gXuVvLqfDp2k1wyVf+5JC+5k0odZgtYRE/w3tl+8s6ak
BiHlqGqyghE5vXeEP9BeDCctgFpmWP16u+XBt7RpYzLEW6v6A2t0qEIhbxiRbK5w44qo0mHJHXn/
VUvvJCuHziQ3/ChVc3q13q+y+CmEM3/BlAmDPvJfh1H4H0NySoTO12husT+7HP0sVOxHzPDQcvl1
v+X3pzACP18Z/YZ5Q01vGdp3nzlHCrsytxvXXn0ih3p396ydS6x3BzcS4Di7Pq3Bn+4ov8W+Sb5S
HmwyfNEN0Mq7ULjCyLJoMG2aLs7005vvM2Q6zB5gCUipQXjgqN8gqSMAfc29AVG+PAlBg7FPpnCb
MbUXyM5a1WJ6O4CCBOpb/1YYL1EiMq357OmKN2wG2xw4625NdQM7Mfrd0GaorAvNm2QXDxpwi1Zb
OwfT5DL21H+wMB7pwBBE3zn0vkh/O5ySMYQ+S0dXEwGeTd7fQaAhGgno4Q/c68Tlb7DkkD/84cei
Q/pGoH/A/OPGWGy8krPGpEUTQzZze1Gb24R/lQe9CZ+GpHZWnbuDCVU0s5LDlraF9zLE4wa9T6Uc
WZyVLuLpyM3tuC3Hf4b7Pk/WsQcVQH6UsrzCe4sPXmIfPyMxy8NZ2vJ1rtBgPmWlj8RpFq2rjXKA
1Qxhz8AY5TW0yk1jAywU65JYxne6E/eNJNGOc6WPBrpzd+g+ZpN79WJIqPyrph4WcjkzKRfgTbaJ
LKzRQ+H3GsRhZU0ll9M8Lf6UaxVqblQ8YY/o73JV7pcnMjNElQEdOvg7wH4AG95DGeGCGSifeQN3
NTJz+QxGjsVggd3l3PAaaHRo+rGB15kSjmv0mAqD6SIW9eACsXczDuE2AQjGGSqESXfiJL/yLzRZ
KYtbMNYb4d61CADf9iHhilXPr2XqxkqgjkFTBxtfYnlrxq9Iq58hpdIQSb70ZYbAKE3X1i2HFqaC
O6QKDzb64NNBrBKS3iPPVhmSD/gdlJG5DNYBFotapmefRKio+ckmJw8HAEYAZj1+lwFN2bD60Pc/
WXUSyju191gDWM9WTe4QTd4YKqMxBNUzq6Smqg0ZXuamQe0ODLAt3GUM5VaZFW+eHKJ9B5zDtzvP
FexxNrxX7V3cbY72G8XwVQrcv59Xa67238JkVok2wk250tTHH3CvS+dpwUNZzxEhTt5MeG8+0eNz
53dXWLR6iiB6q6Ne7z8QAdctebDjHCIAsHw7cV3E8Uk55LTE2dhuUe9znw76VrOMompj5H8SresP
OPn0Y6nGNqWFEXgZKa+NIV2yZ5T619k99QEK0nyxK2ttfAbT18Zh0vpLyyTY8tuz2VB5be90wYwJ
98mVl6A+BOCzNMAVuGvcwlPDZxXxwHmEN67sMBFLd96Wan6QZPYdte2bw35SDiIiM6MIrxU5kjsd
e7znyxLqFbCW+/hitU+xIWL6mV1tklVbzMfXXAt4x0hg6NVtYVNB6xcnElBT33SFFToMUSLp17yh
OPLFg9eo/u//bsTTg9eEP8iK0qfrP9emAdLO1fa3OUq4H9OiHb70pCYwzHq0ku2uDNYBQ3SZCanT
Rhc3h/CRDCcGVrfq2wYJfYy3sHLfbkzcUbfMtqDrwJhH/jKjfYpnGEcjFrnx4huALUQyDQi7MnLu
Huamf1az6KUfom0kp/P9CF5Lox3memhkErWUAW6s1m8Q6asYQMLHUSAkfR5Ts03BYY62VkcA6+Mw
0xDXaGVa3b0q0u0KaVhZZUR+xRkn6mKor17B2bGYcAhRiNJTnZmGPxhJOD9o6Wo2+dFxrZEk507t
Gd6kxfoC/u10GJt1lgj/eBZz92B1HvkE4saSQFwkvnulPbrpKd+uBcZq1IiG4516StBjBpxfRHXY
Qto+wq215K9403D5GK0VhNobSf/CfEebTUxhXTPkuBJcgmUCVkkf+5ONR1/ydUGRjNmv5bQMzQRM
WyeKGmINyEBom8g10M8i8fo1sApA42pSqJgo2RfGeesUOjoiZPdJqpTepzN5MiUIwZJSkwc6uXTt
QALHp+1+QVif1mjObd0jEgrMPkpXBnpCHMvTU8OFyQ6anZ0Fp36RxqkwmLN18MEglne37stTFyJi
T6YK0Wot5fG9XxCRxZdtrcrcW6/G2iTN66u04mzmyuVVoqX6trrq9JjULcZ+akWkUoEshTgvpsqq
GbS2ly8e/OTZJavrDqIc9Yv0/YG/yzsRYdYXVWqmp2DKdt6fzdB6EVLJdiF9Sq8aVxTISUkkQN8F
jNqQTa8dWO3sGyNpcxz+uGQcSwX7XlMDlM9rWF7DKfd9wCnsnqjveXxyJnKV76sob4lx1uBYzNwZ
lPNIZZZ0wd3+odEuqHyxE7U/1kS4dhuS4b5F846/AmBid7vC2/Gc6kGoUwxNrXDp0j6DVEhH3gZz
zhvjnyOyLZ16Y8Awxbrkv/vC4Hsnz2y4HfVtrXfNdUs72OM8po7JCOAamKDLxWhwfySGr6+BS4hP
xLxRsy5lDcAR+7h+k/W51e0OaY09bnJGpEcWyzQLv2GryX1vYF1MNdaUYySJVNlmQ4dYQ89OIbqq
C7JXR2bWzUFEQbYXFWhzrtTVeePOWkb4T3KArBPz+Y4FOq94S+tRxtnQmm4CcPD1Z32K2GVA1hDt
NR4lxpwilPJUs/U29/XyeoCdNA1tRVZrnIlNuWEC7ZF1JtIYH8W7yJqcnEyruE8A2a1zxW//cS0O
kwbxA6a18RjuBUCt7xpHuoRF9n5sZTbQU+Saqep5twl5ba3iuYrN6D0JDI+tmd7aBeg+mLpE2NXP
1C4O/WOyp7oc7+QO/lFwobHKSDY6pGUdq9GfohLO3jbYkBG+RIknLJf5l5YejgiGGbFgC2Z5LYUL
wgoFmb6+3xU/P96uMt88qHZk9GHyolqd1nwOi7Qdmyvb26hitYIf3vfM8UEQKwCcz68F2RRCiAAu
yb4ilTnXcJ5eKqs/6fecDKdssLcpmy5IbS95kUB2JbbJjCAa1CqmuPO7145UN//iSEbH7Hs91QJK
ehClW7Z3fSF2N/SkV64MosSWrffj2p0uoSDPimBT9sy+Hd6q8Si6MtoH/4RFEbdJd6x1NsGT16gE
3AS+zjG+ar/xcJLQ97qaTQ8naYSklkRWjtA8bmVo2Z5w/buijqIGoKpd1b98ImS6b8qpuda7V8yw
+yxz+CRa/ZWE4NsB9p8lo1jIJcd5v6051yYzbQTAmM4DtHqzl5H3rVWyOpJwAUK4mDQ/xxo9ek5C
lxmYacpCg+NIoYse9a2YjECVb/5CeZin+afJpYVxNob9k4jniDjrKmM1nm8Ji0EGV1nfgaSL+FKj
dCfLPBQL/qLuyMOww+bLSKvlAzt7EksMEI+3M/1sBZ7fTSPjyMeAscVAPdZKOKjGc7a5ZO/yaT/F
xq/TOxUW2BUzjRSR1ke/z9LjoT5ZbVu2w9zffx4n8gVZFOJssX/OtDpSoKsDiYqPyUkgisKBtytF
ClYqFxtYNnprIqdGKIffUh0//0wwjjnznbSIYOhJgmDCL+VFjFDfj4UsdbZTKDPX0lnoDE9JlXC0
RYbtZSofLdBCb+dxkty205u8oDMD3OUbVOIVDnuYctwPsphq+3UiuGIehvSoJQ3k9M7A05GVWCFv
OMhaDMA6peXByQiRntV6ygfH8874bhyBfUwVU+P2g8vuMSf8NWgbWDEgOt8eJumghH81SalzN2WD
uV4uHvALPOxXo5n8dUCDPgUqgdeXQWI8elZ2QwEs5+qrdLD7TbiDbrShzMqzPbuo4YbcLY5QIC3E
TjJ4lNZ8Fs7MKN/VXQxb1/3ujPBikjiDLmY30tbiNSmQLf5quc+YjhKzck4XfZPXytOdN/Pt1auh
xnRb+JmNT7Z5ITUB8lHxIHvFf1fOG6qjBHOdq1cl12sdaeX9GRU1f5UYaCxR+/mLgjpDg2N9lH3y
2xTfFVfeMpaAlNUyUzRXyXOOA/zNC+s1QDbq7CGNC22pUzbT7RhI+P59O729gx1NJCJeiLtgxnIa
qoG5I+xgJivzqhfm2/ID5RHaVjyh94/qzVqSXXWV2L+BBoAFQHy+jCoojuKe0SagHJYsIxASE1Ep
72oVv6pK7zO6XIhv8iNsyv28cSO5UCu9MS3dDNX4fP3piwt1ucqOXfDEFBiuT8+1244RniHbRqEn
sJaEpOIk3cHUWGTX0yJAPtEP8241qe0SuBcKgKlQtJKiKdlpXEd5gW+5c+o72aROAXqzF3+8KzxT
wneAxz+Ci4ZMlGrRum/ljXn97WT2i7CdoUn/DT9wNv53BNCEkkL/26x6i6S12PJUaQHYs+ZWOBMU
4ZOUAcz0ASb5PgGa8jPZbaZKTitGJd/spYjTvcllgcarGDm+ZRo+RQ1Pv3Nm+6rbeRooB+pyKG8t
gfW/1RFW10bUy3U/N0+2QNnI2uy9mJe7o65S4Z9aE8IqLIb/qtmNGsLQsdOwGmFn53mC/qqwaq6O
m7K5Bk26a9nDm6huRrI6ju88to8Hgo+Nkd7/h+eVsFUie3AnBBQ4+k/uVEANeZkW/vZbaN+GlSkv
F235TSFN332pMb4M044KsroAcfwIsxIYAmFlr2FdnC98cCBlFhgVMFhGzDnpOzq8pldEZ/P+71+/
RsEyyGrhkfgRMu+lXvaT/T/8vkVn+Pdx6s9xW9jh72Tw+WTi+S/UoMJnrW4jVCiKEZEB5kkZrs53
jxHKq8KbDzDB2tgthYtUjSKWbx/+QxHPO63A+sb+6P5dEtCu2T2+DRacDRwjqPE5YWTyyOQOGnWk
FEj41bSYfv6NF7pVM2rMjqpyHAIjAaXPoVBLO+5cxSXbah3YmgfhX8VaJZ7HPaIQRBTogEIfzJ2W
ZBdiwe0AlIImONEYlQYMaI02ZUElq/e0l22wbwKZY1Amj919SuZXyg5EFMMMbuNJ/IXaTbQkilhd
goltx6Mqi8ioyUdEalpVvgsPJIPviSbmFzJgQ01UHv9seUbkgQCCWXgIoXkIxsQ5frYfrIZyuSas
PHvO70q3nDjtQk922vKIt72AqpRXv8UwV31NDiCdcbSst/dFx0TSdCwuYCvXD218OicEplJtZypS
jH8da+HmEeeEp1y6T4E9wasjwmnfsPsOYI4kxzBYH+rpiBshZ2xF7Z62gceIwcv+I/Q7+TzBmWw1
7CF6BCPW3/CDlaFR4OoGAOkXU9oXjw31HlZvLTzpcFhqh3X4kNk+2lob/tLRWIzp5WCz1GAvDalv
FYgnDf7IbhlYltnkdWAxsJ6ltketrHzOGdqSR0nwHzuolFPQXV6rQWng7Cs2K6tC7KEffSFWs+FC
mD+D7FmwWx1fFMZbHPbdS+745EestWK98XaGBJVyn2qosUbdun7ks6iqKMdA4/VOaC9vqGoNvovf
SQl0VpXYbGi8cOZJm2iEhU1VurTxwBYDuAWdZ8X9szGQVeGcFBR3srKBcUxHCxD+Y0VSzMi4vDxh
TSMKEDY5cJuftGcWqscmDecoyPHS2P8LRwWQnyle8deaNEJLYflMzV60nshpEwD2ms8mkJ/nwDHj
6Zt7X+8DEg2Y25OZ3dQZ4ngnxwmP16++7cmlaB3PDjKEbJL15CIgUeRaL21L+0FeHZbGBkwQYyxB
0fKxzU0n8pEXDDwVC+Vl/b10mSJjIBBJUCI23pkgxTRcNL4beJeKfSc34v93rnvaZgl5pV/5WvF5
RpnWu1N8PLq/vbXOS4a1muGFyXWj1f5IZMErW8SToc3loHnXdSeMFfNRvbv21xm37HwrNE6xFp3n
zVRQizkOYHZnZUGV9ZdeofaAPmYfFA7KAApXt7KXNmxxYWRCvKJY4dDN9WH31TvD2Ymd4jd24yA4
EmozlYerEarCldZJsm0/fnZTg3Sly5aSqBlZaVv/h3q4jHwyktPYL0SgIz1ccTbQKGvhuxkLonv1
i5RfU2+p/R47yq3++QximZrMfyJ3gB08Gks/MXLmLF+Vu683bmi2j+xRMZEQHzXUQ2qd5MXXA/FM
oNbXABCAZX9GZolIJQVj/jQ9PGKN0v/iAlctR1S2ws0+P9hUyVr6zYo5K5BniuUoYljwA5rYlFxS
xS9t9u62DEz+tQJiZsLObyfz4xPpoEqF7gpi9DJmKwtP3xqfjgl8k53Ln357kPJyR+G1xXeRfQPy
bZMOkciPSdSAF37XEWNoBgBlw4ez0EpFEwnrWqGS/puqzyEMjGKflkLmgVY397Y6SZpsSIEhk/K6
2eV43OLCpj26Y01qYS5rFzraPHdkt/MD8bGJD19uDZUI6P+ETPEi7798FuR9HL9WQ5yDOuq7W3hD
IfexiSrX4GmAh7T4a0I2H48aK/+2Nbwis+ChFqIwxnXOO5mEotha4pbKBlLAzph/DiWToyq5BPag
iXRlFT6I8YUP7++Png9Bt73d9myYZ4ozmOMVEBe5wAzbxr649LHRW3wDlJ781FJBk9C8hBtelurD
vWgMgK90a0hyQv9LZOyuxp2ndLVh9mOhHaQ8puUArwTrjs8yhsHnsAjVunTmUFF6Ny8dRYmHhgka
AMc8q7gZm/2kvHxa+wcnjtXsNEM5BEcL1p/SZoBSgAhjDMHLA2RnGtU35P197RoGpwbidMmXwNUN
hj0kLE20P7MnvmnemKWvmwDFSrcxlynkv1MfT0EzyowgNreT/o3E4wNl0jVYsGP6uKRLNEAIUFXV
lW3K32nbCnKcfExqPxFoBQ3z33r1yvkVA4dC76extdinfiJDwpp/eRIqRehW2XL7VZzCG3Jjv1y7
A12SNtwKpxs8+3leVyw2lUhXLz5qr8ftvmOPPmehKeoo/7oo1UxMXJOR+l7LQ/83BLRICK9r+oj/
VFl0a33xik0+2KfqypfWJ/H/KBYCBKdftNjzPdH3fDvSyRmZg12cffcs4q7rRKpKzYkYTrmKlSZy
snkYVyEbkXFFvDqEaSZkoT/3APBP3ZmxQwYOxP9thZURAt77BumSMShMJXnrh09Ec+ATTs0ntoqW
TuXUiH/pldxmOgQ9wZ9+6Gk/X95+n6qy605KU5flXaD1nocYuB0O4b3L/dC8KWfM7B1IcOeuInpV
plUgCAM/yogdr7lpJhjKcGfmvQw40e2ncI+r+9vrKareRcYzFZ47oq115q7vrYL8YyOkoXFQE5/R
ZPpcmjcgWtLwObxh1cJuVjLR+Hbu8QG25l8kZw7kpsiFfq2XNh4PNQU+U16R7mk7jJpI2r8b0NA6
TP59EGWwttOwD8+n4Vf59/Gw9QlSrqUdM4hBsX8bY80Cnk8+sQgAlPSkpkwMjcUZlmdLgnXmd2Wk
VuigeSIn0JGZ/i1YmElKnA4UD0tBlPy/hv09TtJiQ3xAKZOusrbPdbgyjb+SHXc2CHXTde695vXv
wmYSn1Cj6TFsZKrPaPk+BKti4WT2o7OGMO3vgKVFqB832FzRNR19vuPlrt65IPdXBfEwCpC9OHcW
oNGtNczbXNGbvLCvfwxt0sTrn3te/QuuaGXUpZoe9pMXY8VhYqTAHEmbv7kKSac8dUtPzJ5hu6hO
WTPDi7yxloDvosrl6Tz2aCdiyoCBKlzXAv+L9DpXef58zKLc7FvLU/ucVt/925NeEAoKJ3aHk/Md
5LjdaTmfAZfok6C6+J8zJ3DH1WWpN8tLJ/Ry2y9PgiEWrxa2jsqQVSvje9FwiHR9Yv5JskZ0mt6V
DuYlz2SqqF5RQjFHG/JbjxNDg9sTRje8bv1ZG+GaYkIj5ixL7MnxW/CLE2gyR9r3C5IGEZSnVTNt
9YBsfs79jm+dEpAHWnIIMJ4Gtv7tmqeq+9drJW1vJ5IRcUErClpgO44YLJxzRWt1GH6GwtKXRSQV
kRqRoRVCD/l0Ux7ZakfhkU2R+X54pwY6NLuksFJB5g6uFRDChkS1jCvK+ZvWqImTnpxwDs6zro+a
DkBQUfTL7Okjch4146YADL5unHBfDj8cGREapVW/PkR0c91XNp8v8Zp1eNaDmA6YwWKZ6yCh72WV
UtrS4fpEt/Aa+P+nmzGefj4uxgiJ9TsWjGhiuUxqezbzJTk3gcqgkixHLC8DKzYUe3JNaFqGXYmU
sNV2IUWuDOIWkCN851/VRsZOHyVKkmazlnHibsjVR/trbNf0qtnW4UP/QlQ7/1ZCqwXWUKlcbkFE
cIYmgiaaoRjih+yw5lkWyLVxoiw0VJgtM3rlgVg1Lk8h6mLvAjgFF1BvsZpjmo9ikeHcvMIurFjK
+k3gbOQ3NPU390b+Q1HEw/8xcQ+idJNzOhYJaNtnHtJS90IorwE5Xbm2QBnW5TkQ7+Ma4Pts6vZU
rvGzRUqJWzQYzWO/awxdhhO3AHZjSL2paePXie46hcAXqGjp+kLi2B3tYgmYzfgzEdn+TfJR1Ayy
zr+GZqDccVZodQCg4jPcbotUucavsn9uaEp6fbzRTEi7GYAfu1sFuo4AzFfcE8pBQFVIT6D0G24c
nNl+uEw652phDvAHMiPQcVptYXCSllB0SZ0nA5F8n4Z72UpHC/clDuCHgOLwUt8WTREVhZBUpGPv
ftBOe6Si5NFKWCNjDX028XmN3tpmtwYtYwNmZDPTHVETeQz9ROwpmaOQTJ5rlV7tpu1XzzNKeHEg
KmH6hCjgkXHEze/135FKeyl4iTNH7QMdBeOoCwttrZuR8WKFztvQC1ZEqbLLGZ2gT9wfBhwa6So1
PvuvG8Qd2+O8Z+tIdiEF3WissjCrxHq4q0TSPpxdSA8622AVZaxHMj2z5EFcRqxPOQfyHEB9e/dN
q56QIBApuuOg4YL0/65nOqC+f3PWMioeZwn/pHBHg7mN7KrMi8+PEceI/OOGF8hNoMyECKh4Sti9
JeK9T0aRz1KLyMzXgVEl7GeckqGi4Bfux2Hri9BjWYiGb2Inn1F8PcCFESGTJv866SlGe2SjJle2
bu0AEdB2CunveH2GYfcHvG8If+y9Hw3XixK1vUHjaA6KwBf5ob9ShSAL8bxx/BhUtiRPm7Uugn1Z
tLKufdsLgpcTeAS9kYLyg2pMc1nYzg3C1SOjCc1GdsatglCT6ziHlq1kse/JL9+TFrMG6ElI+Dni
dfAvMsKc/bLg55I/39gG8PBaOV+8AymDUMfeS5ZE+Yfa5vPzj6ifmakNlF/ReyGTI8n8UoESUfLY
q/6IsMY/zOvV7J5rmKvV3NsnefetAcRN6IaSUORewXjIjfCv1MWWNJPQdiq9KdIabneyDgubo8J/
VW/bh7+HRQwLQ9rKsD85h8O/F3UMWVLzNazOHfT7M9FTFxwazZskl2zl8AQJcRL3rdUYWgg8Hb2h
luSSbd+Ts9MzEM18uCjk+cKzo95oVxWQxhzDcSR1RqtcXVw4p1TCYBBh0T6jTY1blqFq3XGku+f4
uenDQ1yOcjou324HVyGvjXFtNutVqiufBA5bgAZH7pjjOdJ4vHeJn2lXXo37sVkoUvnQCbG1FCl7
M8Bn6GWoTJfoBKiHMCdtIuwXFNybKvNHL3P54vF1TLqp8Lhfpseeg3Fm4N9VXaNm3MlMUYVDra08
zJMQKxZRV/60PAUkF5SyPj12duTtfQC7FfyqQfrqt8faDaeVEMo4nk0s61Fey3XzL79DYwy9q6Hg
5DTps6aEq7YZtKrJaP2A2ECtu/NNVZp8LHrdN1sdpaI418lW5YYvnVoZzcEKqQgISAgrevoKg7vR
eZhmO7aNs6q2bMycY8Bg9stsu+oPBqm/wBmOFEb1a28Lbl9eLO8qtX0GrXJAQKE/QUM0PNt40uns
2BerI5+y927Q8shm50c5LuPH2/Yg62e5f+VzAOOYurxdnYqeEcnquekBA3SD52B6ytIkMP8+Wf+r
uTrN/xyILnBOmNDEUxiixYYSK8s+9p7WBbWW4oXvuYfEKTGUttJIrOaTqsb132Unyvqf7R1YzDZc
GAwAA+JIQGDEqbDYm+0dZExEAk9tDDYcX3+fGMs1MQtSt49M1auSCNiT0mUtVNmEsVC+nVttPXld
bxiK8Gx5M/sL6Qb66YXj19RJETtZPAP/ffQ/o5QioCtt1LXmTDMbcAp9oM24mwrYR58R3DB0tF80
bYbvA+bhAchlpv0b52p0qKZmywugHzZYo1L9Spr8I3f5ggVutuse2f4YasbszJXfI5EIWMojPnqY
34HeoUUd3pA23DC/lqNEKVs6F50vW1Q3gXEVkudWGLefJ+e5AvBDIbOtKgw7LrxQSsMRCoyeWoKb
YN97wdl8BjxnMhI5j1qZEKxEZFA7b2sKBpgE+mjfTjfNh3UO66S8K7mupIhFV4sT4pDz5M44LbT6
bmR7w9ygAMEgs19JcNPv3F8vxctBzzSsjszjYU+74s5JJKLLLRDBDlMzgA7gQ+v2yryiQgI20H5z
8172Y/971nUYprZAAAPLc2HfhbywAdNyGaHOIaAkol/o6/r8Vt0O+VM2kct/wtexbxG973DeTVU8
1VnmlM4RGiSy9nCOxXmGo88VHzb8D8ygQq6oUVBIsFoWFEg7IdgmbeaB88Uv2SYWTpven2wULfYM
G7H1hS4K317GPbCucBNqSH+OvyEzQfMtFR14uJM/TXCZ6oD3/5j4YYbZC1x/2SfFpyqWMDo3hypL
Zm+f+CSr8hmm/34EohbkZvgAGYB3xHFi7IG0e758hsDZp9B9gr1eYSqZ2PQ7nn+0FOEy+BOgnnTP
mVEXNis0wL1enwb5Am2gwyO3gBndkicwLYf7xgkkRk0Gu6Zv7TRd+ctlof5PxAKuQMzXkDCZZcRf
FBeTZlktXmEJfKTVLTnzagxqmnfQd/mnm3yOdT1+oPO05nENatksi7fGV/MbjW+ovP85yUbrM7lF
bHPMQR6DDtWo6DF3O7DpeeqG56ih0y6VvbgyJ5BvAkWKlDXHS+HzThoNp0KiaVqYqNvDep/S7JAM
CQSJQRESSkNCJXuDrHmWTMmEBvjCzQEN/L2j55E6+sofgHkOaETbb5395I4D03FFHho9qNzWRLmj
w+3LN18jIhvRY6JNdkYyaz3ewbrXU1h2StqZfAottClL/io9p/b2O1mGqEebOm7HyGQS53prr4F0
lD6iLg8TL8xo82isVD1UGeNxWI/dTQUWOpdlIPdqkQBfI+iM23W8zYwDa84YvU6VEnGbj+RYxdm+
+fTrxKfJ8jmodeJlCSLKcbMjUZhAUr1kRard3l1OjhSzUTlyzdyvMAPIAWL8ZmcV8NhUpZs7sC1Q
XejhcCoQY68hAzrjer7A+1Wt/z7uMnvtENJRVAeBQWfj7BLQhSnwFaD5xPyo8pN0WxTTBJ2DsWRw
i6VGGlv2axdZPiIS33MoIL6Y2ocfyNidS/4BKHQxeznW0HYWkLYyW/wCrcOLApJCIU4UZ2i5YDgB
7ntaYtSU4Jw9a7cypHeYB/eZ1fB2HU93o1ZF41nEx9a43qasWETSTQrGD1J+EpqRX1Aj+6EEZRfc
EbV5PHZJ4PlOKMOBxU5dRK4uauUsCpp+k+AXl97QsAfQ4IOf+za5xMdozAJSTsG+cLRmaO4FEsxW
UrUysdNgs9LHZZbJsQMVB1UwLDKsK2TEHj06AGtpSiUMeEm8pXSDXwQdC6xZJtpvLVkxc+P+eou2
X4XNDFpWAN9ni6cdjhL/Af7P1Fxq6rz0PcvsxWxNPjaV6ecQ7KMGhZzwmMNgrbx8WteVy7/bC51i
d8g7Bvv6wA97+6zbZHsIVOLVfnjLXPzRcdepUL1t+LXb+ULzHwFvSYTbt/1QjkUi/s7PsJPCUHWC
/79ImXZ31S7Odm9A7dOhImgKLhbkMHgqV/sKEQLosvfT5rmqWitmICT0lmlEpq4zM/MiAfak59md
E94FoL+KF61eJ0AJX+z/jF4+8KwtjPTDI9hRHy1P65qRbSogX/mFlXClke9mFHmWHcDP8IbFVCuy
coiIDIy15XjSHn9WTjniUkWfwQ7kTXLPlOvU0pVCWlrqTzET8CVHbe65nT7dE/a01gQVauHcz3PR
y+Ad42QQwVsByDMPY4es7S+qd4sMlMADcpslW+OYL+E9CyPuAukUyVka1WIlsU0gln5988a52sj+
skHJMDV5ThHULV9J5wF0rpNsboAmVtWBX3566uZVZtEQcheN2bt8czrAluQvTnM5MDlO0PTiUxCr
C8H7GrOwTkp6J/KxSvSrDDGeXGOWc8ACTprjVYinD1neLgYShPeHqmxpaGTE6/irfZqGucQGXqql
QptK++k8kiHVaGymy8O6TCJnO7OyfSv0JIB5PpOUxxw4obYKLIi0HNCtLRKIPLQwCfQ2Q0IZDiZK
5yWaKNmDQcb2kGNOvafXSioGawwwVg11QUEohVowvP1hZ1BHQqO0MOLx+Y33TfkIQPHi5eGL7dgd
bhkW4tz2Stmitq/gSLF+W0RH5huit1Nxj/L73Ds/cpUE9KxZfqyTH51WOibiNUo55CYCZbntcEuK
q7ey6tN7XXqE42j9MvkBovm8JGSdeaN1/pzbxFQZRp401Q0NE6DCjiLDai6YeO/hPy7bXnENJ3tA
MDmmdMD47mZhfOGOdrOvGN7xbtYwRHHQBIa28FfQtg822LEXRH7t8ShEqnoNDjerLeJd93gNihwH
Y+v5/tnMFChIk3VKJn5vP3DllYBm8iM5xIvvpUXehGnJnSnWYXyrfq6/8EKJh1eF7sVxOtM6fXlT
KsXZI1ptGbXYyGkn9M5cfA+0TwZ6rwYbGtDroUnTPxZy/lJK1dSJ44VIAIbmhjzXFQdBLXQzbqhZ
OE79xOz7CxSrOW+N+E2XbKrjHPvTrPhhlWKry0UBSl4EmpTolgRCJIquXYDjbeBVD548fHNfLtNU
vYDQknyimNFcVRppttQ2jPxBTFgaqE500t/VKOl8HXywoXjEOIJly3Lnrj1Urcdch/WgetkGz0LN
SRyHU/8wTwJC93j4a0Aay2ewGVBdaRbH6ZEOaqPSQlBzPm7Bdg5MJe2an/lEe4VwKWLxyNfFaHZI
MkSlq9IrswTvoKK4G1xzUkCMO2sWHubaOY5uXxiTHXu3N0fQ50apFfemIhUK7iqopoiuUOrPv02m
Cd1ZfysY6HcRDKL+9p0+o4teimexJdgCj42EaDquQkT0C9k0Ed9tFJezmxs1VgG/1R5CD8CugfmK
scMwoSL4kIq3NNq+LXMPiNdguyAUb8x4j3X+JlI9yGCHGFHW02WZ1VQW4tMqMjO7MRjQQPRZPt7z
3taQNeattky4t6X/5wmAuKm3E/Tj6AptWI6gAkgUG3573Wj9w9+lt6pzvRbfgY+1VvQV7nf+XXlg
E2vmDo7h2CK7B2ppMYt4LTlx3Tal9XOhEmJ4JL0SQ/vv9pGFwu+CWD36rz3nmBfBVG1Hu+kuAobb
1XxBBL9O9P/0AOSm2EPhQCR0SHZkCh33zIr26RAHre3wIDF4KGqa3KHPD42s5MQQ1ymbo5YMxuj9
VMBRws4l3I4tHxhIv1+EL6f7Xkijd85lCS4oiXema9ObEH66jTkj0nt/62+ITWucjaJ4sJMiqlq3
zK3fIyidPEv8+3c0GgGuQl8kLvll5DxhsU11YCt7R9y7d2Es5N5CUW0mpvmtk96UPfzPoRjNlUkz
mLP5gsbPBpOul6jjPHg24xGvGF+H/a8vqsWW7ETI8XUMxgnyZs9xRfKTawmoj1XG/flNDj5YDQJN
9iQZndoh+2atwp/BqR8gTlZ9HPQTqPfvSUISgdZ9Rr6L/juiOUQtjwHpjtNAA+oDU6CSN/G9bhxW
OWLOXba5tXQwxrLf9hS1ApK554NJqKlQF05CMJU75y1kzBEGiW3UyVx9N3tqbtiNmrnujEHF0XAU
XxGTrBh8FHgzXYDQHGaDJWWQimU+qm6vYvhz3653ff+VBsmisOn1obnYogGVM4Nw816tsKGT20ND
HGGN+qK0tjP+9ITElQ3h63zjAfuPUCV5c9sp/64QV9YHBfJGB71w6KJbBeSP3cbUGrG6mXfEVIFH
tm9zIkYikoS8Hb+GYtfXlgEaZsvpjl29SblDrNZjtF62EfPp/Fb4px1+VadP+up9GfkWgOWv4tbC
ilOsFt9Vabl3EQlAm1kMsk2dNDyplsKaryPlAWavsfL/ooWNK4RvsGGjRKtOU4nbaAys+eLYFYMi
niywIL0JHmOfZO4lAPrEoaLKmzE7IWy9CkVxCkRsE+pORsATJ7CGjyPnCAp6ooT2W3IR0tOmN25z
+v5A429zPZrmO45gAeS+YQFlBTtyLCP2dVehEAzLvaXY1ARnG+Jw4t5GUEOP1rkUtDnzhNiwl2PV
Tt+h9BZaNu8wM6Y9FkiIQXcx88prj1wU6FeVHR69KRZFhPogKu6xTADlSfJaPMcEz+tvboBWYkPv
a4l6IwUNqEZSBab/8SmhDLDgjKqQcgGMC6dDKpKCgRauXVnDqBNlyGcJjWDUd4ekChESsQoNWUqK
qkgaRT3dxhkrzgw7nCwgFUAxq9hS4HCgr4bSGWza3lRYlUSdiLXj1HL4hJi8BsHLNbvd/s47uP9c
QA9jONbX48Ej05IR65lsfvthI9fDH4RZ6r6aWo8lES9hvolj8Mvhu7/YdGzpjVv5WJdAjwL6+JIX
x48YSdWSZeVWqr3Y2Kk8to1vAoVN7aq3FEnEbkqeVzdcAiU3+gzjb8+/qEAnCoePEv1gZ95/n+KD
+UJL9/A2YMj6Vqdy/nUOiWMQFIU3F6I2LD9TqShv56e3XwLJssetw6NcLznysczdbpJFXVT94bCT
8YjZuxkPAXE2aRh/X5FCob3ga4tg3Mwc3asr/Yuchk6OKq77vCB+F3EQRnG4YbDnaw9Un7kGipHE
DD8MCbp9zU91Jzy+zJkNU3KmdIszH42I84lzP5x4Hcb2TAdEnVhZfjjAo8wr9SPxQe5686CqEmvX
9jsaMuNNI8/CnxxnK7OKB/tK1yQPO+Np/tylhlVwbX8x3alxET/dNYFrVRs/CsDNjqYIUP8kbSkC
75gDKBZzUPr3tiybgjW6ZqO9JY+vLJEH6NAPDT9nzKDim1TRHkgdzPxFjWfbCIVKWSx1LwZvFvxx
VAMU48ZA12Gug2v65iR+xWYJzofXLipGeoJ875nIx6f52Pp3/NTgJ84PllGUZcTd5spGqkf87hze
dLTAI541WM0dA2dPhjBlrw+tHWMASlTc2KfqrJ0pfCiRmW3ryk/xNva6B7Co1HQd9rw3Vtm4vOVt
sMiQlV4ewHPJip/LKg/2ZGx6xrOkCszPPVSlNfr4r9pQYkbru0Yl2RizudTg+CEcdq+yjjNRyf27
9fxuRsGGuckpEXwyyCXfognGPSoSsBx1XtEOG/v4izCBhzgDzKplKYli6xRWQLdzkEv+9w9j3Kph
roRUMbxj7GvLOniLh03i/yY0PGye/0xoxgz0AV8aI6FpRxIXcpuP8BVlFpeQj2PPq5JPCdVPr0KQ
OYvHV/YzKkNMsnCTXiqXhGQfrlZw1uPnV1PYgJsP/SIePBFHHQmB0aVYQ+l2IKozIcv/UaemtwCl
AIKWH1c/Bl9I/tl+qsjaeu2yoKRabGVSSDKlHACMOI2VOCeuwfeFvz+CMKqQkGQqcYrVuU1U8hmX
LNenOTGoS7p+ijyr5ZO1nAcnqZPbKBi1qV+mG2fysM5oObIJdR24cVx7eXvetaBI5nZMlwoZD4Qq
jA8t8uFvY7t6azgxYzmdSjTdwzqEHipG1t2O+6U8ZMtoeX9Yb1NdIRW3SYsv9xK63COC/RNwdLt3
iLrxuAqQbSLr6wGSYjNwDc5VftLV7Ruola+SHPtNd3QsRb3ClSQPCNU/5O9dKzNYKB2dkcfhx9jM
LGIL74I1TS3l2Rsu5/KnWZOSMZKlOut5nNdjzoeyeay2oWRjaNDpZdpcOk3tMNHa/ZURrijeFEmY
JgzGRcXsp8DJTvfMmziujG8EnxMVHwoC4SakIAB1tqfJTuyYJu9VjxjwY7Y5Nkj4SAFhyDstkfCg
XMoCqaSTjwdyHzqTieTuCAduW29mHbEn5dgcEgyv3WKHtNZ/hchIC4m7kzoqcGF7OQwYl4hUrN6b
7jPWhfUsMR3pyJlTdnuTfI52A1XRDIut0dUyaFBr3OoReCtuahFiLhG2gVowwzG4TyPBF/8BMn6u
iJWpE/6kdzs7VlD9rFAdeciBRdrv/cl+cDnm8rttdqPrsamwgk2knbp/Vb8yFNVJ7oGmUahc8T2M
XgoPckspbY3fBXQ1o4Li7syAeLny20VbluT6jUwEs8ZnCW4+Z3q1wMhwWoZ59VNUZFt+NHYJTwlD
MvL+O4WfXcOTlqOy+TZU27RTtmXANkQVz7FeTTLJvOiwy1fq9qE4l7QZNhTR5kYPVcQE4cE6qba0
EiocJ4UVZYaEVxR62nKlkQYESm2iK+ilxCSPHbPELMuYws/6W9TrnFCnO9/JysGn/XUAyHGw5hXV
cS07lmjtYFScU+joMaeKYfBXfTwQ2XCC3rlCM4/2eO9Q4Dalx0BDzHosO3lBGF2LEPD/HsqRV1ng
kElDEMLDbItZ97hw6opLqfCFdWr8VupuhiZ/1Wmv1T7itoidWN87oRlNV1sCQ26QR4Zp/P39K9Mt
XE6UXivHsylgQZ6/Vi1TEQBNyJvynn/51xNGOjfCGlZbkrq3AXdF/7maUUiprtfYkx/AF9YgZqDk
wKCI/5OOvujGqRqqi8N7cDhDhDlbo3CRB7hWmNanESYd9fuugjeq55ZgNxVNZHOsvi9Dtefb1JlL
zg5rNUeheNR94tw7fN0vqC2WY9xueGau0GyUj/D9yRLXWP9cID1EO7mLq5qwEKX1qKeOR3SjL4dN
GSPgKliA/OHDvhPGeha3qfeXJ8ZqZLP6oDmrIS6BqwQ2PE1OUdRrmsL6B2tqvSrKVKn4PMW+rYaz
jwm/Ew5Wt4Nng6NepVkBckJ+DggVRU8ajt9sk482eYbnqEKDka9FuDOosgeIri918MNQXgQyRXGo
P/Q/jx9ROaBI6c7bLFAwEPTBIOdRjuwJmHBU0hfJ+fcFSkMU9ULvnTTJuhMvv0cku2Bb/xqlewOK
H/fN3bdCAuG+zyuIWMhe11ZhDGRXhbQF+/UaothUBve2nMqzX/MwFoN2WV6l6SYIEw1HWrRHKcRA
mwcLJjUXoT3tEK3EqbTcSVo9N/1TUcReKdXVNRWiBu6zhnff9Kz4Y5XhqthnzbGczNjBA1gFz+FG
jlktc44gBWuJWIRZjOcfIrUNCkv96vEKFTRoAGJtDqcGtEHo48DeXmA35W4IjatWfN27Q/nvstyl
nYgfef8OnVE0FgRIU9fI823gsPcqoH40VU+ua6cWw54lABCkqDomc0ekxLs0BG3/nKAUW1tt8IQT
h/ch9seYQz2842UAXDholRn/33uSY0RCGCLCPpq3irKlJQKMk5aJ7Eu+MVoVoiw/ju9GvKSgA279
wzkeWrf/eFZ5S2Iwmn9byj9SGfC5dWBkgwI4NExu7qUMniDJ1jRKe/k0vxLNGJ3+L0bSgkVVQ0Ku
CMbq1U73y8SXD22E/QEdNfHrx6AztMQkp4vVxwlbLintr7tN08IeFNRd3pSwkeyMyiEVfHgt2wLk
2AaYvkz5YyLGDP8PsQp3blFZFKYgLCeSphgkRBz8H2SF0IzVL8LrM0Bioo+3tjpZN/iyKv9/R0iy
zYFeNAIOI4qjK7vTPGI7LWCU8OdU5rGXJdxY0/CUidSf5owpfmuMLhN3IX/kSITumA3Hf6zwfDT2
rJrxDktLklLxqnidJNPGYFcAbbixPMe4a/Irpfba74wrxt+UscwJixpceCP8eqQlHDVC0sxtMKpi
q+MRDJuTL7+tbNCTFrm2u4InbnkROa/WRO7m30Ct0M+W004y9yRi+JsxHUwUblfDs1xtTd2TDm6r
bM4/GTVM0dHQEGblQGr0jTZOvMrE44zge0o2dXJXySzH+qkDk1PM5efFbXTc4PNZqLX0SuioClDZ
hS6iRNk7KBjbslJqCWWiWzqrH9PECww9kjCMrto5jxHasXPHG3ikXwIQCWmC3FCl6uCzBQphr+mw
hQtx2HM94DlTsuige2sMmwiaOAj9So7n5ODWZmjoc3r4LxWxf9aZD4qieH8zg2B+d+hN1Ha5p/4P
P4PzAIFh6AEayU2YZir9kwW0CMur5R9fsvch8zFePGpqDfNq8ybyGsrN8jvJ7aMdDxxyjhdGhc3z
Qv+fUk5lmQk2hLZall+LNqLEf8RV8SV3XGZgP8vzYJqGXhZnM3gHMtpDZd2S2qCgriYniwxDzHAA
rWTW4SHKgJq7xFy8aKWFAuqDIrn6x4AsgCRaysnw27IkwgniWCu7qJI54tbPP1MlnIhezjCSJd/S
mU/HZeWZKO1IpkXSPkYJhnwh1scij3zYZaOo1n4Fd0ZiOPvm1pDWYc/RqsjRXnZyzdowT25VFoZY
gDcjG5A2yO7e7FVNgwnsvx9Wousd/5pQaq0j2TNwqz5TBDc6BPZQTRk5faSR8PvVZE8tpmAkHi2H
3MfnC1YQpKybVIa0pQPu+o2XmFmEKD4F6YPOqWCQmEKYjADPf0OyFPMHeNrCaidPb5P3RDXsnpmw
XM2giJFk9n7FyZL/slWEEQLYPfnGc/CDZhyJJREnDnh67BREvv6ocQ5nv7ezw2TciAJsE9BUovbb
JPkTS5/yBxrs9kWdEFMMqxG/bb6PWg/tTwGiyc4j2yPdqvItW/gHRNELo4XVgdEbr2TDkC+NWR6a
bH7LJc4pPWme3c2Zmujl948H1CokwvlDNljFJiGjOt7kz4HwNFiwWNrhfys1Gwk5Ay+fy0I9yZJq
Pa+XoOplEeqXeVNX4xNpu0LXa8IG3a5G8FLb8jXbfucCsX+kRX/i8OvT44W+Zn3pNHUbKemqTQZR
PwvwngWuLvleZapAWVB4PTs+Jm9QuD5bYRZAAdyYwIpWm7I6h7/7XhyEB7tTzSkAo6TkVR9DCNpi
q7w2DwhfyuajX3FL/iUEKD8deQ6rf1BIJ6uIz9GnLJTtzYO86DYAE0T7xzncXEcWoJi79Z+tV3kU
q8hphvXUV2GieTGX/WycYDvm48743mk8DDinuMkpL0oWuxJs+pj4hLw6rdM2ESJBK8L5BazOIAG2
02ejb7Iv21bjp91aP1JM6/XIRzDi61KXt1k7cA1bsZMM7NSt1jAz52Wqu+DKzs3OeWzRiuj7SA0Y
Sd3YmHOPGphoIhuIEm4ssThUBUoxb+IyedjoDeow4u8medkvigkSxznLNaAyy+lFZUpYhZfA85Pn
hf3KZ7++PTWecUNn6n68iQD6CQIsZDkVnyIlrs51p510OVKJDv1UZ9/mhIVwBHTIogy8ub1tBDvc
XMXg32eFlR543HSnZmisXJi36MB9g9SGz++dRA3NHh6/75NcQcSzn2u3lrbY3vDy00Rw3gEftTbe
IfYM3xAwnkPVdHoDjYmKpDdon6D55dWhGZoNra7MVeNgWAi0BvOhOKNemG6h9huXUcN9a5Nro9Bu
VvU1K6uJFQ6Ifa0U5qhJqjnk4Vi+6oMLpPxy4BtAvKM1tOtldgwiqTYIYYYhAa0q2VZbNJDQQNUX
jjQVqRLvyASfycMXnqsXrQR+ygFAtaIBC6X24T2jB3V/ZWZDwhGAZ0egNd7NPf8+xWEZviijsyqE
/4lmMCKx3hJdsP7ad7lMdAnXJm1MSzb9IJSxQAeEnQHip6nm8NjJEozMK0LdisdjyyW8Lb8rMSad
mtesNTNard9sVa9WkRPDl6dlOLZoN2GhLfgJb1SkvMjR8SF+d/FATibyswbNBYUK2YRkGMd7OFVO
i8MuV6CLbc9Dh+yb3o3uv2gGrFFGqHvKtX8UmvjZczTj/uXzkYw9szImdgfXKHgc2MnbtLcyCcgJ
VONzRb4563XYWoREnzKynJL2qAVZS9hmYrlB5HIK6vr1tGtzqeAM3afaDBjo2kPDOWkDJONRDHBn
UcuWC4aTHGASVsOGWCOkDzovtkTEzB+OLrqi3H+7DpVRIMlPqz/8C/Gzc9K0R4uUZE0eElHB89F/
N1qeXT/KlsE+hCsdu0ZlIJapzYHhuJ2yHORidMkXlxOUj4MyGqLX4U2ppzTIz2B0HQOhkO9VSrLp
MuIwFZB30i6Yy/CW9qvJIcjOTYtQu4k2cGuSnkFOHnHwJiosElC85aSFsaGFbqwo4H/runmD73TO
0yLy8uyIZEekII3afIW+g/PtsLhTLHPOsQX5jeOkwP6BWqdwjT4T88hzjoQz80LTNDOITijbf05l
dWTc90+EiAKi+1ITnTBnhrF9Q1dcYLsO6AP812yjBfViBpG+t2rh5oRcOQ36Lr9KFeAQBUwDZ2SE
YPeBJFSICKGaeuM3r1ZsW6AEzyzmK0qzKHis8kmWSf0Z1x8+RpHmlTlplCEUqqNhedIPVi/+WAUJ
T2w17xioy7YsNoPLF/x1xjuNZWTAizPT0LvLZkIDo5j5N+rW1l9QaVj/V7SJCAEStGL8O8fGTreF
s7e5uDv/o+tHZMqpt1BLknnr6yGtOeWl2j+9QHeYJOhjtS62tEg8mKRaFWAbjfZ7DpgCz9a9Exx/
h2rhqGmQEVvoO9ZR0jAGuxqmLnnLkutvw75UxOoYbokJHO6dh/5UuivWgNfbc9AI8FSUtIN6lv9H
c5+l70196v3eCYxRx6Z3RxxEkuzSweZH7jgCNbQjyciLOvUmADYutWtrrChpqwKXx77H/dric7Sg
Fq1h4ncJW6BDU/1SmoPfxLX5vSOnvBjmb+IbkNUUe3mfjbc2OhTn2A6MbwivFdmbZyaxVIAwFXp4
8gEjjWW4jtPsBR/k8Nir1/BYu2jjEEadHMKDDScU+VnMwIl3yXTxiVmWbFkGQoFA5RIJjEJm414m
CkIjoCU8aA9Z+pz8uHXI8K4u40UUw1xCY10CMIzv+5GAzgt4THN310GSrbTUQudB7d6LORCglvpB
5esE3wrlsdLuF1G4kJeHUj/4fnyNJxLQveHJDpfK3hJ+QyFLuBzjU+uM2ot5wLHlieyev5mJNHlS
jehrCzja3ihgfa5i/hJ/V4hVGZx/Exbz0w1rfaBXZtrWD/Ml32poGDXGEQyR3MAforkR9auSVszG
RmV8kf7arkJAIfR/G952kHIEyQxHQJSWHh7plRR6OZCCTGm4rBCHYYuP6cRuVmtjMx6KyyTJpZVo
ZsXiEIm/GHVuTngGYYEXMDnB7hhxnBDbuo6FBZA2PgymEK0m2vvJsjOzJi4wyVrqgxMB5fqshsuD
w0yRLm6R62lhSweOTLYFJ/ZI9b6UUxFP8mQxDRqZSamwzSiszKe6ftJNJa4hyvnB22bvyuFSH5Yx
j+1IjYZr6evVUyDlsMMeEmDUI6FEeYxZSPPfhm6lFtjWQy1j3ZojToiV9xkSAVFcVRf41fiqR4v8
dhvETkExTVg29fZjlvykHapvfeRXOR2SlyXMcsiXQLZRrLcFg8t+uaMs7S/El/s5oTdz9IRunauS
ny1msDoQwXCISzl5VBEzqpTLovbmuAaid8uh4ZIiGxrmN37VgvjUOVPVCdOnUmJDuN5wnzWOgcVy
vRhORbwc/91EhBPjxavuQRCYVeBTvRvAvYv32XO+7F5hjNtWTwXK7gUEXRshwN7LhfGkOpytF2k+
nOvrQAqc3CRsqgiR4Ye0Q/jdcIFSqfk1XZOZCQysApGWBeFLBKJMKbKmPLIzlS1DAxp2RVZYNKry
C13Y6a0WN2NKEbCePgWQtN28osTm1z+6OFUZ/GVnCmHI9t7bgnLuG5LiFLy9w8ZV8n7vfW9MxNSO
OkPDH36SuTx924xNALyy8KCNfTv8qjxMeZGA5AcF7u9uJgzEVTY77CBraoVZ5Lva1CfrASTRW29s
VbOGlyQ7t6TXxnNq9cpmPOgvsCB3OABnpiBWgqPWWOMTDMzn+bOhK2DBPSVXaxABqskL8orrDegd
fcUOsUjDhkshwd0WVqnKU82vAwUHj1XH9mytZSMoYpe8sv2Bb+8M7peBgTnd/nyCF6cSC6VlTlHh
M/dj1YXPEsxO/L/a5b2uoTqbU+KwA4gyFHvayrXLR1XDxwqj8ojdLbxZCDNMPWzvWz6kSrz8yh7m
fh64gmlJRu5zaPAaFyZeH/slE28laWoO6Og8CdgpGSdRGAIrtSd5rlk2OOVQN1oy2SLzIMKMJG9G
kliY0S8e8GcGKkiUMmC/0Lr7BM3h6peZzbjLTVCBEdvTN1cqn4tPjwiR0iocRy1J5FXQ+/RtB/gZ
E8UI2WFC1Gyrx3a7lG9RTo8vlzeuILyjz8MLoygn6tWUPStk49xYAAc/YueDWb3O3fo+8vh8kdip
VlVJU5ldON5FBGRh+LN7I13akkWR5ElFPrSvPbfWgCLCubXR72NfPhqgOPWcHxdhhtmTBtCdGCkP
oCoPNmK08CblezNPVvkl9h8wZWBwO5TNRENnJKGYUZI0SRKvEcK+W/YDgIhaB5gOyvD+TWN7fR6y
x6BzZPqJGzBm1KgOlFO5YcF33sxpwXvwvnk+vg/0JP9oOGuE23nSCDHD6yTmVAkY+LhDmtjFfhJq
9wcje3OZn7xzgspYPjbUF0GceKg2CDqbuDtIJkW1eDpno5A+X/3nunt+vpZByFQ01ZYPcPpXmeg3
E6SascBQySAOGaM7YFr0oSzxJabCd+Xu8QoBMzsnBwjg4/pKZPTFDx7kt6le7Eiiuf1DslhZ/OQV
eRFSBB01S2/6zb46Es42r4POAxqRvDyCJ/CFHVIICNIrr9/jpSLNj/FQ6CQnhNhI5hjPoe1mdlF8
qKXjWnOykeRvWHePHpzu/ZmBouszI0cKwrwf0uH7u8YJIi0FhBJjOnPcs79ebBTZkJzCLZsql0aE
vEj95CFtx++wzCiY0JhnC+g001rRJuuXeWofmv+/zeGOFWgyH5OySZ0139bjxZ7g61eEOu2N68p1
wJZbDHbXqNeX0QlEByEOfkT6NRX5Vm34OrbVIH/321SxV3gpXqk6x2O5u5BI4jzneZ1RIXvxC0LS
vQfNAUk7G4Kuk49ILLUTTmDdOEg357CCTuuM8KRaLHRd7s82hQaUYSQXV70jpbWgCXmv416B/gNL
3RptRcf+sNmFXBG90D9xFbod+c4WUoNit4LZSYH9TTOHs/t5g7xxA7lcr9oNA3+nUcbQzVtzV6HH
uly86eONJ1tCRFFW493jTxtEXnhQ0RPy4GO5fwbCWAKF9tfyaOcqyoOSW2Zxn3CGd/N3434gWPpd
G2Ev+x4/lPUGs92TZs3s9T3MXWJScQRgZICLwhDqEChWD0cnpE5SFo56cmFj3T7tN8TIzlRAqWtG
cpQ7qhLC2bd1FTebI++VUKsAHzegGwLg54KwotnN2g5DB8Xex2PW9/H8am5QAS5ZJFmXX3TqX79K
qw34i+k8uPuPxJZnUi/44gQtJHCX9ae6uo8ywhCbNN0Jg+in/LF9nRcz+nRdWyxaBXo+YKIaZXin
H2R2CHLP/nENK1O3XGhA9u2R4c6CzTEMNIbr12jOm91UCWXrgd+oNcq6ucleWRx3cCLJwzpi5JC+
Ey+d+eqWsjMAl0meuYEg8I67bdJ/rbqVK0Mf1iOAWkJpwfXHMMcUeGc9IjTYRNmhhtnCPWqTpw7+
MMlBvxTGsz1rnSxJRjHnLzNiU4zEN3UZaEbcjrAtrGxCBpv9fGCaPtdnZgCFZsbA9i4epXxJVDhy
zIP9UMrvMjglcWpXS0pA12wU/SG+2yIGDfWQ7lw68H3VHPKnzffe1g8Aygz2E0QlcqIOHLt4tTIb
Vxyzf7Mvyqe1pW3cp6VlN3bi9jcv8CGmJA+6ebmBTJprOw8kCR5qBul8L9KGOENPF4b9r3WekVZc
Xx9hgo40p3tJVGWI34LY+AI9Pocz0aX/hsO+ZqVN8kL9BZlm3eiLBR7p2Ew6ILggoycqeiYHDyFf
EWquxk8UpE84R6v7jed5f6iPtUrm7dlrIsC0ulZd1AXZxCcSxF7KWWEfCngyLAa2A0QwmLb5wuhE
p7bTcwhyQJaWVL/m2vmwzaeiBnwmbABQpAEuSYU6/sjvA3fxjhGOG08YnpIMbjwf+TMCFpvJpJ/V
sEtwZpjlg+ssTh3jcQ/WFEEtbkL/xfNtkvHR7Qe8QvNogi8F/IRpSwR7tzqzS1RGU7mu9ZYPplCg
fRUvQMFzT5TYmWEgKxzjyg/UsYKII8A1PnBLv0XQbQF3DiT2j0zPr1zVPYbkY2q+zEFshhUog42X
bxZKhc5ggj7vpZbLmis9hOo7jzC4uuE3PQDwQ0VRKYKX9yncbPqi0SMF2ajswqOxcEqcLWxlSQ85
O6+8kRkgzlIRehonfsCJNr1PpniSDZIrG+H8XNWaMNsqo32I/c7K4eHmfHjZGXVlAe+7Cc/zxa/B
IZt2fs5Ejld/Jkv2NpFglUq9T3YOmBALgJZRgyQhG0f1McpvbUbJKxdqEVAYkuMQU2RmbOqHP9af
0/6XTFsPPpE3UZA2iVAJdClKPINXVWbYslfNuM3fctEu4vxgfcOovUoqFgPn8Trh+6h8ppR9v4Hi
u9zzzt/T3K9JzgxZDq5hIJSKhYQzGXyhaN3PSGK1/At1hChZg6bzb418/WC8ZanQRv4Tdd1d5fFq
gKEpv4gjD+uILL1veW1cdrJzKXbSkQPXE4rmz6rBAGr3kmHioJAN4DlhlXioace2QmW+G6p1lkAJ
mz0QsYU3pFwpHmnaptrfJjq3uIIIyd7UmQCZ22lE8yd19moDmcNJFFLF7BuGFl8dS23QDhbXwqOa
j1ChNFPHjRU47ww6dDEJFydMFOwpLGgagEnlsgWwYpyym4+UGfIf2ZK82F7NJ+//pOUN7ayO7+UD
UWsONvpUSCoHghJTQmeKM/MghHXXFsWvOnfiTfTrOXFusMiTxXODI/tIMFLKwH3v48IpnpDxKXzc
k2vr2JBGI/VdwPoC3fKtijQKabmue4DPgg3xkVraIzotqJ5WBk5/Nw6ZqYNw1g8bvtVY1nRQnQw0
i/tKNbduwx24xnOG+BcJ3Fb0tO1Q+BTlc7e0FvKuTceF+Wd5p0J3m56RNMm5i2YIMM8OT8wHtKRr
Fp8kUxpKSXcuUzRXwpJECmmdbnioWMK+5ZvlLc2hVbQgAzHXZ2tgfoWI77x3Apr1Iz/QOQzgDbKU
aFUFdQYfCYsZ60887XjRxGUOCutJGfAfIXvVtnJAu131dpHQTyXmtoFK6yONuICK/oRYd/Y/nxDj
brqJ+ynxweoxC/BB3LvaCFRoy0R54QgbBKdKvWDZNTEXfjLF+3ORPLkWROlSzhIjkJWpkd2IgSsa
ytL0Zu+SYNBERzjUYQGlTOPubRXf9CB7Tl6PLY9uq0Bjzz0UfBBMEKGsCBhn0y2WdWsKcu5DNSwh
7/G8UmTw/1jwG1FTCugQ57Ar3tzT85rkZFuDi/qg1GqILG4AZSqi74jzp6whNtPJzCgD50N8FrnD
p8ycxdDLsGIhvnRCBfVlt/Voej7wGGmDJ+aaIpWyA2g8PWlVBHY08dhFoSQAnl6SloFgz5Z8UE7s
I2pEJW7S25mNwQ87KtwCcy6ZeIyuvlscrIOTuUxwoBGob1m2DbnvHm8e5dqKws1ecpyBsNBMwK6m
b5grGASAKivwFiVm9LseIqf7cQi65k/OVgFVBNfQQ7fP1Tkazfjx07eUhGBSYJyVn9HnbDYeGbvT
Vv2xzFpXdlttHx5Q6gXaL/teNyuFd42wNFMm1g21iiTncljVvwd3XtXfO0YHi5ts1jxIdQeiqT4w
mvKXb3W7a6h7X9XC/I//A3NY+2Rmek93JT0LUzu80i6udnQ43aVAXqBTSycJTWEswWRMJaCLnapc
LK3H3K4hvtWG1CJS6T9qbaCfjAEdm7wP4MwfJw8AfgxMGuzxbncVk5YEBMMfKYNkYaS6CQ9JFkxN
XqVga7vX6D9aOl4zNPlj7Vpc88/f5DKdjZQOtncW1szQy/ZVUGzT1W+wqE+tezTVg8FrAjpPIvQJ
QBjX6z3b03ooKFhRg4kQAEgkiEvAsxZ+slIELLhk+sCDLqw6Ir5Hiksy2NhA+HV2H6Z4gqUGGMXn
195ZqKDMRDOIVVNHuN4EqZJav4+iA5nDVVTjPdJn1sYBCvt25Fag680QE7gQGoGirzy7w/3Rych6
dtznPNKsLEWLN8tt6mx3trpUgTIjNAwPXynu8KferXf5OZMS6hjZ/aWQtLtIw/GO1qoadJQCQtBA
aghGZdm9aXX/VcWyepXCGVbxkcbkONnKJ65iarT9Z6HmGOdTEBMtWB+TC+0FlTxLTChczSh9kfVJ
GxMQD/1W81STk9S+K6TR7oAYsjEXbWybzcceY5zxtou1C/awVKvG9Qbe/ykxHkpjsDFcIu5wo9On
clnFZ3oI/+K+9vh8gri1HSInkp6dKuVocrKeVBRWp9xYRpFETOVJc5e3dL/85csM8KeuQRN6LLxg
drYt9g2GxAGOl21+G7h6FEdfZPlY2ZOjKM9+V/Rjj347QluWc3v16tGrf2ko0M/k0TPwQSXrtujC
TlVVupk47lE+2mzPX4uxf+1hfRvXwL+QBkaLbLUvkbxDlEGFpTZixgzkipZq5G77/Z+tnWmavCRj
Fj6HkroAfojmRL4o9qYlu/yD/5zwXafGZwhnbq/Q2XiQMSLAu4r5m/UL7Lq7BZxQIfyzLFpul9Ea
w2VAioDXiQAMN0DHn+DNOl2qgJKO1VFf5eQsQDmKlMHAKs4x6v5fHFjzTqq3I93eMZh1c1d3o3Jj
LelQCYY4p17LLoTJRibAR1TPdn3Bl3NKxeT8nq/RB5kalSKliESTnnV9h73MrypAfHx6gicpVPOa
ZFhrJ8xzZi0EnWoDbPvzlDSvoMKak7h3+lTqNST4XPfjy8ApH4SjhkbkHv/5C+Aa0GAmn+2osm57
zU4qlD2qe1mCZXZ7ZyrD/whqV0APD9gwPoFY/0/xb5l2gEyXA1/0fqWtcHrLKKhvvKm/fz96DZ6y
ae3qZ0EqZFLujGHuvro0SFVmrfTeA1c6mQC0gSqhi95SHalYodWgUl4ZYmwOACQzRk1TR1bYDnsh
WcSoyLWUqux+WhfrUnSmE3JPcqWmO4nkrHHvpihGYxWJjMh+lWGbg+ebUN14dHmjxuPMQJri9WmF
Rbp1r6xfLtNtiuU2mVhmVjWZPf+tBWItENmqnmMOtvbPqHPSDQr1q0+lZNcebMJcbo+aClQZEYPi
+0oFtqer51MsjdJKdT0iEz2eEjjQwZ3O7sDjzzS75/PxxDIibi7I2oVZpukNJW50MktckxbdFjtc
yJPbyJM7oLhwi4srWVRWK3E2MPjPh/0mgkiQ8kic4OA3+sLw4Q8Iqg4o6DatP0/v5DH9qUlJbr5x
wZfpBZ07+xXXRHEBeAMMmuUIaGAL+c3yWHbYCxsrbUudPiw1KhCGfqjFxtxzywv3pKUt+iZUzFF3
kUjmVZA+I59J55E9QlDeDZvdeSXMckkMUxUzlTS5ZDFIIRQeBv4HRazTFkwCDF2dyVbqC+oXijMB
RGu/OVjZwGogrVkJEb7HxRC2n9V9L74pkW3wUY+k8+kLaGDTPApMuproGju1MiAJJYIXIBVe+GCw
A3mJ7S9ZZkZu0srMbg6A6UA99wi8vDQX1npFmlXMifGBlw761GkSJevc+I9l/W2+2zId5XQCvTbn
jaJSHbkN5d+mWw1Gufy6XfCyHP2MA2aFj+8NPEB2XqUdpRVrp16ZINbpafwV6N5CQqXAISgC8Ep8
2rCSTVvNgUKmgU6YS69l5Wzo/YdocYoJNd3Aio3NyBD4H/kXDIbtfElVfv/VQ2v+I5KdGC4Rrtyp
lF6kd92YtW2NUTC11sHL0yU6aIiAaNpcjGKHPJB1Rzx6hO/FO/mLZ5WjXQV17aTsyjEgSHXtDiIH
qrsvLFW7NH4W+tDRdE45ZhLpRFyzpTTAMrMxr0C/LbzgEPqH+2fGYAyGWa2D+5SixskenyDNJsTu
hGQa2VVMyFaWnke/xW2zLpMrOT+eB3Gp6fMBS3PWzvB+XEt84JGmKmZiDkOLYux4Td6EyrfVctCN
oNVLaqWeARa4O06JxiPSgXDiPe5dbuR9ag2nZJpUJFt4Rr6S6YGzCwamJKM6C9S90HOo/Z6iCaR1
cEw3UsKmtu3wTvDix76G0JSHF7YFDqmZM5++Ysxy8Jk9K8dHbbfJpSRuGtPfHsNIaAbUAaibSqMe
TUuzzy3YyjtH16EGds/yY7OSwAYozcPDdoyHtsnZV8xphEeLtBCyPLEPyd5r8n/klmGtxGkaD3FM
47IOArAuPmqBBL+Hdg1xwmK+IjBrIhKKbg1RRsVA441tV8A7BXpF7a57buHwBgRw7S0XgZ67w6fW
iYxcaZIxhwddcPspRo3W195BRuPKMOErR/mU8zK7lA1sXzvfdskNfig3JuFziW+rOJJ6D3/qH9+Z
fnXQmd39kca03OuRzQKwmKXD/0aytLbHxhXJkPEshEXWAOvgUIWFAIE3cYzWUPyS4Wu743N0Zf/p
jilRcJaOlfU1lwmN4/5sRL1QG9TcdZ7Roe+sD3Cx6ucTmy9RdhBk3DGFHT7sVW6gJV8C1OMQ+Npv
1QbuFrBEpUg/7AmnRLAZWjIPTHcRMJ6kSZheosLsW6pO9zbxwg8PWDngq8Wf56kdKF1t9OFUBEjn
ESICUh4fhqz1V39eb2v8iOTpNOe3lBUXpfRnrf2aV59oM60MK9L6lwZ3zy+oBnpqGMcupQHVF685
0Z99tCCbF7F8qZUFc2n2ITCzsCKnJHe9qehIjDVRfd0HQz2mqLDP9h1SBz51KJMr9mE1sg8kEtQc
XE3aE7yB7lg14ZurRGNex8V6XyB0tgiNVSFeha8vzwAJ745jRDydvCezLueEE5rCsERoLRfrDhv0
IES5uMQ4HTHLe5t5PH51ZZEdhwopL9Evh+YmD8/8h4C0VKqA47FUZ3uCBovNkfzAeTYfJ2eqQdiC
nV9tJLikr4j07GBQwoljlVFIc4E+5XjFfaEzxWPG32NlymdnckZ6r5sN05FpfLJBEqYu6axFTjrd
RfTvVtkxruZJFgCxkHGbyhoRJSWn1uzpP0HkA+BY8q9oqy4695PJkwm3RTra+FXcI7VXjl9bHpwk
HXvvqFy/d8MWsLL9HPrCeSMslA/8cMhG2SFpQiFzZL9a39aFCZuh5lAJeWgY3Jqtjle8fPLX9pMy
ToYJwToVwq0pzJ0XtJqXTYmETRRpGsQTsU+5dELIzGTfwvatZuenpdKAP+Vq31TAbMYSqjmMs0Sq
Q33k9OPIsEgTk1/cIiZ5ldSZJnbVWBk7nIWhvUhYd90s15TvjZXAZB94dJoxzvHjIBCHApjhGzoS
MUtrVFgurjMuE0T5V383GfXNhvRuXKA3VWAm7Mq0ceZD64X0mVCAYloWTLtC9Gn/o152zlDbkWVO
mhN4UV10PIzVZ05ADduPzJafWkLHJSuVm2u9CQUgeoWCTAjvNSV5MZTVDrXVFhMkQe3IYmdpuDcP
rRQ4pUFhIdnqeNOEJ8Mbs8vtN14jdVoUvMZ9fU89Lx80KO8DBW5pT0YKGR04odliXm5P3UVo2581
Fmjy2WigJRLXJQN9WSJLpJkIgauQuhMacgjV0m3QvMvYzNwIBTogdBDNbKmNxM+SVm+JhvBr9/Ej
QppZyxIRmxHe7UTyPxMgOiC+o8lf0mNyC3/+YlFgHphGoyfY+sohDtOFN59NF8dM5dAduIwJrwXU
bQM+bsPe/uhsBT+bEn14IRoClL+t4cYCWNwnALoI/6IaQJJuHz4DE6bA4TwRri6NTkxuXZ6JAhKn
zfbpBkZuO8K4PDa7c0BHi59hlK0pFruN08DWcAiMfIcANx3RqMVcnX272KYP1lXYhGmPlGk9TDu7
sBkSAwPbomxt21HxNm0lb5EkGmk+3VdMSXwOVDdwWqewMedWCvlX1pOd/ocUMVZpsmF8mWFexxvb
AkBhVGPAbdS4Gybj9cZRYdbHyZKEtpYabCIeh60szSafb7s3Sy0Uil0hntj/yP2FuX3FchRPZ8QM
DoHmAd/eTUFj+XZQrO1FJewAaqNSnMrwxWR0DRrgNOnBHqenvW4jbPn+IMd3J0s3bJwFkFA10FfY
yJq2RGO6OUNz5/rY//VbC1V8Gs8OG8yl2u3ZZPigjGp57J4xdy2BjDGpRV0v4ECU3ycPDatMygA8
LErsOyJEtNhKBX+ZOxYAzhFJojt/r9Wg9V30hMORbBY9/WGdiy4f9E+rokQ4W7zYplanEv+6/lyo
7Bv5oUDOAqNJx6arFPQZNV6TKMLc9HHpE1uwIEzzBnep4yok5GfXbRNLdJVF0SaH145xlGz2dvto
9zi/lotxe+jU2r/jEQTwr9HAGEFCGaym3cX0eYXwJYJfyzaWMPJXj9Ts0Eg830xYq14lP+ODSfrB
ccZmTiac9+thyQ33nkP4B7gBQIkFL0ks2Lg5xv01TV/4jK7dfih2VJWaRLUTIac+veBqgwaCxn43
nreuHrUYuElsBaEgJJUNo2RvANSRWo+ZP3xcG5yDsvaEY0Dxr6uBkdkj6lbqBMtr7jVH5+N46NjU
FDwI7cas0ZpStvvI5vcoDLLAMTERK94pCKGmpMBM7AqtzIxIU0g9QDs1ZFkBah7zlOR899824WPg
9i0fFxQuPorHBY38YsN5MLQvUb68Zt2K1OHvG++Ht2kbJ2T0uTDM0n2vIc9VqwWCCEnCnsIRsZ+e
XM2d3bYqOM9FWxPrnL97cSlQCxuKMxtWb0Of8Q0gNnGCQX4bIO0UdtdkDDLox9jKt+tfn2U8RWL+
BqckI6dkh5cXa7LO6HdtH+L6MCBw9UcZI2D4hgj8GpZBDhRP7cVzLmEz7qEV7eZygpi5qK0rDttt
bf5f9Yq+ygsdglfPcTc3ZutM6S4MHZHmToTbUVq21aRTGXcc5fzKIA/I9+qA56Ylav44GnEKU6z8
I9thzvd2ONPI4iD833s8YXxfK1SWmYfdOYXmiQIUfumCaWqDDFicY7unwtKHaqqbUZpOXmz0Ve9c
//ISeIMWoaKPh//GRu1XYI2hvySLMoBxZ3lewlebTe8gQTvKCzVoOzoIg8bgsoHFMCg9QlOGaaQp
p4hOgaCNItbd3bt+HAHFH1wjMw8qvDE1BuUz6eUZ7/u7Zrs+Dc8szcnHsq059V8tplgU22fqSxvX
yHDxm7Ue3FlUGEZ1OY6JZerJPUx8l9lU5eEiEtEVzhQxfX5tmwpQEmmIHVuG0f81UrOTy8RbPBDA
ymoNW8k0KETXuK8Xcvnek1ZJ2NGGPKUDHI6w6sa7DBofBJTLWlPdETs24kmvxQGxv/ODJC7WHbqA
njjFgTfdPecd7cWsEwD/oNFl68LpZ9x9Ld84GXZRr4GeGu7Yn6CxK0x+e2Eg3cU2Q8SYXUdjqOrs
0owiwxBC4Z4C/piuL5L/aWx0xXR6d/RZnpmcd5YRmGGwJMOOlfSZeeXS2gAVfhXlENNuFjnznwpN
d52/cpo7MMVOjJP096J5LPRuRnaK0YphxLz9hh0ewjQVJJ3DinRJbEZo9KtVLLFRm9mqHzDmytIx
AoFPs13P3VxL5Xry5bf1AaiFtgyoYlzg7Pjs4xIPf3xcTwIpKB5jPZX78DbqkYWwGuHPJ660Tttj
xR5ohJkfr9XD5SMSXkS9u+1GtYGEPO7Q6fObJM0RPCEo3DwqnhgnWBjfHDHm8ERcuODMew1J1AgA
lKxh6uCsKuC6AWHXA9n1VNDRjA6lrXODqKKK9mMddKsgJEUrUzLew44Q1pzmOTbe7nDqvEoyQ96K
vilip3cdTNQTbOpmV7+nt/lGdO0u8F/5dngbYL2zlftzm2M1Wp89w5XeD7AQoqCraOhPe6nh2XVF
o0dNrjM/7eFdEPpi2g28K7Jjv0zEj5Z5caLOkBfnfHH7ozq4mYGvDuWVE+TRdehp6PLkxkQBIlVC
VaGq/fDo6THvZ77ZlPnmd/HoDZtmAPSq5MTiQLK4hDOy/vOeEwaT+SYahEuLvUasPSyWfxzxQM5R
DDIdp9Xbs1xv8in9TMLj+feCXPCwZtgJYwI8IjtKtV5a0VAOKnvYOBlrvRh2E6TBop+IExekw5Cx
u+YDoXfDpyS+gS5VKU9Me03MJ9MOGrhaG3XDTOETKIBLCrjJ0Lclz6zGyc1HHnGX/bt4D98NT6Qm
V8I7ToO6aZCGSSiF0b5v36E7vu2lRzOCsATNIekQ8VwAPJHpfDWQnS/8RsYaVxi4lq+7jMHNkskz
F7qamSxjH6VHGCi4N2hXvt3BZ0pgocXBepk7wMurufKvNZ99sd8xBs1DStWve0IcuzWsEeYSMLPU
DWSn3mc05LDenbSzXVrCtVxLRBYmQFxvEoKdIsdiuhGyoMcoiiTx9iaJ5/RoUzU7aj+1ERyuNECr
HuvQ8j20rszrObVWXeHd+zXi6Ec/M0ZOvBlOhEZVzadk7rNZQuYXmaQg2KrDR2/uQGXLgzRDm2F8
dXTtT3aUWpb3VnxgrlVx4Cz1z2mD9UbGEH3M7IOY3bAWgQogutMqC+4mGBtdLFcFxoLUNbvgzk8p
XuK/M+H8a5jbm+Qf/bBMKzAd9ucckRF4CHzRk7Sz0e048TsxQZ1f3A/Ap3EmRYmnFsap2U6W9vAZ
G7NwP2QeQABZ0I8sGjSCn0i77UKMG9vfinoe8JaF06DDh5mZLndzSmxGsxSVYarT36NMavO3+HLV
9vmeyCrOcG+dzNeS3q/f8vsnaRn8Ajm8gd42RgG0vHZ/5RLySeF8LbI9iz6zc0Iwtse2Y5hy31Q8
UO2jy+qq3KBJLv/nPB1cRJMrqj1wuRBa8yoT9WrSVWU070nK6opSS2fef/hqhj6xupY2Ix2HvB+y
jezegeLBL6r7Kg0WP3k7cSU51EGADFbTK51QspRAno0SNFCtlQOgcvRdDE6/sK+sTKc9JwU+Rkrk
90reyJqwqSx+C9OW7gw6vj/Oaa1RvxduQL6Fybu/a8+Z3DFfG9KLt2ls1tKlfyOuCtMnYjIC8DM3
UP3+mbySdyev3RoDD6ouNM7epg0JYXHgiBdYr6LZoa0UBwiEj8qaeE0qyyHpHGuUBuMCigcK+Amp
mSpXKWdT6Smtvrnrft3HIeCDfe26qGRI7LO2auGXIlfpjPqq7H60QlJxmtYInWjT8T2693+9U6m6
bejN3A8jBxGWcWlq
`pragma protect end_protected
