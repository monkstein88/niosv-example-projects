��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���~�`���sB�G����f�Y�k����f�N,�ې!��
0%�I+���-5Ey9����K��
w�@���	G��"�QDlܬܼc}��Dh�����	m�p�+�#�����
�zt���_��u����K����Fﴘ'�}m�����;��A��x�P��p��A�ְ!���)�L��kcIߙ%;0ƹgס�S�0���ռa�hH�G��]S0!ɦ���Շ4��8m��k�9��@� |�ш��hިt�*�v��sW"��\����;�����#ey?)|�,�W�I;�;B����T.�	7O,�7������/�M��T�A��>��:�j�6DW5r�
7��؇|S�+~�,,#z�ێAAi8��m�|˗`3w��/���ݦ5�I�ͺ�Wd;�#w�Q�z
Fx�����0�]��=7�J:�iQ���5�A6Zc��W����e�MI������sK_��C(����{(�
Z�V��+[ШI�f�o�<�L��ֱH�4��`�u��53'f���
,�.׌��ځ��X�WH��`��#h�������[
��E�ȆN��(2 MIı*wp�@#N1�zjA .���GW���o�aϨ7�[a�Cf�=Q[�D���08t��l�mƾ�1|6�u�@���ϩ��~��^��aI��&3��Q �^P�c�ʂ�s��e"HמAY�>�3=3�L*1(O<�����m
,������|,�|#pD�����%\��)r%�	̈�2FB��b�(��%�=sOe=+���ڔ��q�E~{X�y6���������^�-Fu9Z���#�)v�I�]#Atڠ��������s�j��~�4�X=�����<?�g�q,����I����Ϝp.�U+��l�ƽ�H��̃���E)�;���C{����
�]A�3*%�7'�x)�rSHZ�K�֢Y�߾6P�h����	�é�C���=C�����gy�7;�z�b)^�S|�:���0��j�ȓ��yhj���f�;�PMo}�ߚ�)��t��*��
2	�[Qb?�'��2$+�����C��h�\�~--��[�JW�3�(�5��vÍ��s	�T��0��_��!i9K��e�^,�Ղ��Ē�k*ӥ�^4W7eL�$�����i�J�%��:�r~���e](�[ �F�[���*-.�Z�N��fZ�B7�9�W-��NGm^�)R�_9%_^>nW�b�:SUi9aGɷ@�s��&��Y`6T�l*�|�w�w�"�>��K��u�dN�j_�=.[_��K�>�$$\�B{Iޥ�i�yRtAɌ�1ߩ$�q��QaJ�Ί���ho�һ�c������(킷�4Y��I�%c��i�eq"h���8>�����:�u%���us��n4����G	���k�y��K|=>L(�MЧL2l�@���u�
uHN\S�'��4�}�tW�j�#N�W��@r��?7�����}�p� �mqO��V��u��b���% �L�a��:�$�WˠEҝ�b�O4A+�vR��e���6}J~��Ib��1�o\�����;)���1PlɓA�Ϩm�z��lx�{�C®fY�~P˫ �D6a�XS�F~u�&%Y"�����
�3do���!���z׈2�����_d���@��n;(���gWC"}Ϋ���0�4�����x;��;4�~�KiZ�ܦ�Bp)�c�X����4!F�`b]Г���,�=`\ǁ�+�Í�9f!1e��z�21��h�\�$v�Z^C�P�V(�2���G�t(�Bi5C�����hsk��ܤL3��)����;�GI@��j���r���5;m���	�9��?GX6����X�7%����6��L���:	�[�('�;r�z�dwK�Bw�:]�-F�n�|b�%��C��_i�����⩼aI�Tz�is!jÑT�b�ԍ{.g�L��aQ?�z �*�|��L�ޗ�cq.+7���3A��D��,x�yO̱-���M�3T�~��B����Zv�Fpxc�9_)2NڮǓ56_P+�u�UG>{�sj�y����0�_�����y	�j����o�mO�9���_K��y`���pzE̎ώ����٪���������;]��j
}pi�8_*c�N�s��y�%y�l)�-p��3�v�Ex����c��xҳ��Y��8��n0Q^[�|.'&� �9�Y�2�4��,F3^^�k$|JK����^d����Y|���^�VK��O�z�IC[:�'vQoRr]E_�BgRlw[��s?�h�<�h*x�#��R��p�>��z �Bi��[@�pͤ ݏs���@Ag� �s<��K�8��#�4���a�2��!��KP��Jq�r){�Y����b��Q=���C�����oj��aԱJE����z�kY�&k���O��ሓѽ��.��~ه|�OGA&-8�<�&N�}��#�E��k�w�m�C��O����_���I/M���hl� ������5d�V���CD�u�ep̫"yOC�g�?��|F;�)P�8�����Ɨx�Mau	�m�9�X��<@/d�qo�/Md���Q�s�t���Y1Ԩ$m��Le�����9���J�3�o]K'b_���R��)�_��w�u�3�)F��P����!�(�T��Q���A�݄��~��6��<tY�31<#42��؇r!S�ү�s���͔�?	���YS��^�k����C�cZMA���BGS����ж���#��b?1~~�N*�K�د�O�G���u��QyY�14��y
f~��x;4�^�G���8#8g՘k�W1O�cn-��b�<v�P<=H�#P��o-L�ܽ�^i��"/[�
!b�9%���!���t��u�{���|���x���]Y���B