��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2i�>�|�"���K�W2��;#��Q�Wa�["�����wvbe��#%��ѯ��n�@�"%��}�+�M�JǄ�� ���,+'V{R��l����x�U���Ea��A}	!���7TW��z:�ROΥ��i$����B�`�+�i�&���,�Bˀ�[��9 ��d��a�1�z	�9�x�@�Z�
o��R^y��6XP���`&�p�K6��?c�]H�g<Zx%;LR|�Y2�U2o��:��0�*Lîӷ�$n�����A�U[����
�_6?�^)#��Q2)�o��������"3&�Q�Ĥ9A��/������Ll�����8����8��:�DԾ����i^G�T�R�D~�e4�Wsf\��(���IM�?X ��!e��p�r8+4Gz�m৹�bkF����j��>ŵ���MyM�C��A<��3�1�斑�x<&$�����ƧI�Ǧp�1�ɲ���CӓǶ�'�*�1�[`�ص,ʈn��s�{/�.`̡�l���0+�Gh�DcK���AՃ���Xm�����m4�^����;s�tU��Y��5�~�,,؄L�}\��_
��p

�E��^��l=!{�A�?�<��7�݁�V�5VZ���j]_���U駿�Źn��r�ĔhKk-4�T���]Zx��*��l%i�n��R���>��S�h`�B3f�m
hL�I����2�i�-DF��#¿4��&�p��Hg@j_Q_�{X���-
�iص;�>�q��Tm�Tvʖ���I���%u~dB	<��Ʋ{��b��"�(G3Bݪ��k�(�k����}4�"/��8�֝F��:-��;.�l%���[f
ê�Jh�x���d���j��oN��q;�μ�2�r<�~2@��Wo	=��f�b�>�)Y-%�(�>�;,I0�S�� �d>�_N�R���6���X@�#�d,R��ĵ݆24_r9��sH�d�-�\7���O��sr>F{�ƈ��t/��X�$Fl�*��l�$��9
;�ce�`��I}M�O�ٛk{�`G���O����aY!"ˈ1�_[.��&B��'��󺒚��~�|��t��)����������q+�f����2�S�1�N����g����6$a���U:e�<��c�܍�NU��#�,DN����>]�+'#5��s�*�%i;ZI=Ŧ�0�>.U�}�j�?�?<H�N����BҔS�JTo�F<�xk��t*�$��ө�Z��6����A�8���W���q��٩��ӥ�h?��@������������6�c���]�ˊx���[Opw�5j��F��T�\X�Ŗ޺����.`��{��*��*ݜft�F�}��̘�pi���}魸�(�fO����~���K=`V����QRBl0�)¸�9޺!%��'�b���,:��r��<��D�r�L�"��K��4QP`[`Pe�QP�}w�Td�I���`]k���h��WmR���,P���w��0�9�((*ο��s�1�ذ��g�e��J�C{m��*X]9�8(1�+��"E�M3�'%ÿ�;r7��0^�:d�Sd6��а�pk{ņ��	��'�>&�k�E4uq.{�\�F��2�Ә[���d|��p�ћHk%��'�}⻔��6���b���1�f���ƥ����BT����va�zT��<#�$���}ui�-�Mu� z)���,�ؐ�����; Zmn�z���Σ�G��ڄN�R�I���@��'�?�|�K�c>�)��?�Uv1�k;��8\>t	8�U?��0z��WD��q�٤=Qg�&�.��-�����#�F���r�;�Q(h�oJ�q�K����eN��}�;i��Fp6g�v�c�(ŧt�6wu���a3�'���Ԯ$��;��6�CG5���k����y�Gv��X��C��Ծ��;�2#n52�����:Y�!�p��w�i}^f^vNֲ<'tyPJ�#�1&�~�Yʟ1�j���Xsr�u!@��;m�!� ��=�|�",��laS��dݜ�����3�!(�6���b�S���Mł5�$�;�.3� ��\E<k6�,5y��S~�R}���:��F}�a�Ir	��_�>_A�Һ~�s�I8���7����r^*��l'S\��2�5������K}��OCEa���W �p�6)D�`�q�x~��R
_(y4�nz	Z�O��""`le�C<�=����=�8��I��i���Ce���Yt���f\3�iV���.�iCLR	A&�a'�򕚸~��~��d�Z�f�>���s��(w�����D����\���@�B�jF��hr�!k2�zFU��Cre��F�=uA��ʳՠ�~��g��%\a�i��o)V�TR�c�X�����w9��b7;B:��M�����C��ۗx����
y(XR<��������kiL�����Cpe����nn���A�7+<�2����ym���ux�`��ю�	�]�s��^�yU+�M�%�At�
m��/<�Q�.;�m����"$�̆����!\ܿ�b� F�߂-a�+R	g�I��o�h���vA���m1$śQ�p��o�̐�2���,�����.7Lk�������mq��2�	�#��풧:L֠Nſ�{��Ga }.���0�JPf��ĸp��N�ѲI]Z ��ġ���%$I�F5H%���1s���%�qM�a��}�i��]���W?��ϗ�(��Je:l㭦Ӳu���99q:������H����� rY6��o���&���h�]ec�9��xTE��@�ܮ滻[t�U
"�z��
�6��2�����A�w��<
o�q����3v�<�j��1-�IrM�Z��+"�A~�5�LG�8�`ҙ��5j��yX*����D�P�n�[��A��Q��O ��ZO�լA�D%jR�Y��
�>���;	џ���b�L}rgq���8s�V��5��5��B4wb@�tթ�
��%1���!8�0�Q�L�|'�:T'�6����]GM�ξ<��A�	/���_B�5;������gp��	�!��f=�|�{y�3����㖩/�h�\���l�Ԥ���v	d��>\�n��Q��(�L�vv����iHt>�ZX��6y�	�q�)N�@���|�����;�����w� %"Cs���\m/`GtQf <j���(�Qם^������2�l�<
-���p����.�������n6���?pܘ�'sJ�|�p�"�\�;5o�W�/����E�ɶ�*⥈�u~	<*��Pi�w9��w�/�`9�#'�s]�:�c�D���/U�R�+>�>&/���e#���c���
  ,�_E(w9�i�2 Mu�V�����&\�a������-{ ;���d�x�!-TX��t,g�6����y$��~N�g�<I�
A$	��B@s��؜�ܕ�h���sv`-OG��J�|�aW���t���;��"3���V
�����_d �z3=i�d�x�CsV�G��d*��O�c�+Y�PBy��
?
oRo9Ul�Ö�HH��藫��tE»L���H�5ޯ�Qأ���VL"G��;�� ��?�'�GV#K�8?z�W�fc��Zc�����;�ҭ�f����|/��s�j��=N��L�6|�LjM轐��Yr���DR�d��N%�=�  ��Y&�&���]<�X1�DݤLT�Bcp��iGF��0 G�#m�"�ea���Y�y�TT�7�[�C<��E�f_�5�'��oA��Ʈ{hP�4E�M9�j��_�AM@�Ls����Fv��l��\*�?�L2G��%~�|��,	K��F�����KwR�B���z��[��P�RÝ?~cX�$02�c<v�_���	y�vD��P�M	���cT��D����+qۘK.k�{	~,6�
;�T�q�:�G�O{�y����������{bt��ds<�v������L�/StL����w�ʀ��%M�ُ�5+�.jV��zf�G#�Ne��[#
�u()^h��+�����Vqx�\�x�%Զ�$��˚�޲�����g�m�YAyp�Ig������(FY�0]��{,WU�F��W�������?��X,�e81��c(!D-(t�C��3W�Cr���@�twk���dǂ�������WO럣�H���0:}�Q��\�~sn��T�s���$�$�vB� �Vi2`ޖ�d�#��M��*�UM:��6��ş�8ݙW��%��v�)B� ���ť��L����pǠS�M�t��UC%�����;���X7�	���x�Ú�wh��6�vy,�+
� E�t75����u~��v��L���u�R\%�Z^n_�X[*eرČ�h�<�Y4zP� �/���n�1hY��
+Ĝ��f�S%-�2=��>���Qh�N�3�?�!�q��R^�Q���g��Q�L��F�}�Gֆ�A��D�l�4׉2�BtOU�o$) ��d1���ވ�w�� ��^2+�� :�Z	�x�ȹvе�Vm�U��L��څ����_�w�\Bf�Sza�����X�l����%�1vSo��`��S�wʚ���{h"�\{�1"(*��b勰�_P��)@�A1[�0j*���}�f�s����I��
>Yf)(����黙��=�����㬌�W����u�#�nqi�R�U�������U3���!?���&�!6���Z�V�f̷v �4��k'����B������� #c輑韪&����rZ��ʂ�B�Wf%}�7�3c�\�(}�=�@��aM�_!?\�.u�>�iP�("�/O��3�C�-�Q����!CQ�س�1���捚��� ��-!A}���`J%&W$���.�Fk Q -d,�(#Jjs�P��AK�Z�W'S����u��1fMJ?���&9���.K'��@%~�� �`�SS-�h�����&/(�O*��|��}�EW����V�@��m���v�38*ѝk;���5y������"{���j5;��7��@	��Wz���r��`,��c��G��*f+����*�<��Ba2������6�	k�}��MTw���(��;#A_.�(M���	���(�ZP��U�>?oK������iQT�U�����:�"�ԋ����i@r��Q :W�d����D�M�Q��W&X-Қ� �U{1H�y�w�"��4雷�Z�ȫ���ьT���
���#�Wq�����7��/L���C��V#�_���-{D°�I��⚟��ʾ#��!v��4
.����F�+8�@qm�gպd�u�l�CvD��pk7`ǻ���$y3V�|�;^*U�=�QT),ty�-�� ��_�*|�����fa2��ک�O@C�'Ϣ4<nEh��I�0b"�ߝs0�Hf�R�/)�ӫ��ݦ7��M��%x��C�w\�$Vܖ��_���7�{��\��r�^�bnJ�� é��)r�й�,~���	{�{�)���^Q�G�6z�u�jn_�=�A�.����|��T�B;X¬D�"#ºz��R(�.���dn�#�w�6��G�e�_@�Y�u�uyTJ��0�oHOf��
z����N�	T�mf�-1�@Ŝ'p_��؞5y��e=P>S����Z3��j�N��ZC�� ����e�[A�^�K�����d'��0��G1c��^�NS@ir�?�kY���)����bR�
.(�}�`1	��_{TG�g�s�E��\�ua����ԸA$E`3��\�����$�'�u�Py��l
���\�[�[^��ӿ�o�`���v��ח|�4�D �� '«��r�c����dy�F\e7����v��]��vn�x3inO5���	����������)����%y�R=h��ıeY�۸a�}A�+1S�6ƌ/���B��L�F