// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
QgcY2+lCPdQk4YyO/7tvKJv5ehAkr0dgCbP4k06baAZU/KwpH0gEE318peu/UZR9k5DTRlZP/2RG
Nj4iG9KjZPXe7CIYlVTql2/D5fKuoAffNUi1FiYyDC/p1JXuPEay5LlpyIvH4vtx6ijI314j8R1l
TptadmNsChb21diMiaEe108p7R7XFhk2MyGCikjF0yYpt2ROGZ2LmTExDIwXOr6mYHS64W6pLPrt
lCH6g8sVSoWjAxodKD1/myHahTmlAL7vbo5n68B44rKzO6GekBuPmJOFyBQ4DwHeTikRRFsbnbBe
xzSFNG3qkV9rbJ2dQh+b5PbqwBMz7nujjQmMuA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2160)
dbF0XWLDVgjSJbtNpG1N59HQ/lFYfSsPLwkBEqztW56rTs/V6MpJYxtBEkXGMcJ2UHUmp+8fJRfq
a1PKGGVgIW8EqyLXJub4NinjiK9shf2L81GMi+gZprEQDIO3jgfEmaSO/AUn5Wo3lNovzLEq4030
heu0+v4lvr6SbPLsaM9VKR3DeeGBA0t/ldE0AhaGxWpxC/qvsr7mHJcAGFUbzNrKnsByASulLtsF
atJurkwqYP3ZDXIHddJ4y1k2aKwwoT4kELc4zudVZsYtzLyZbQBm0kI1X9XjkiPQRdtS2/1wInfc
IogsClU0viExDmLXHkGk/y8F4LDiN5r/H4wcruzQhiEQkuodok7pYY3Ni3G0hAC8vmG0IlN0XI8T
fcx00VwXSF8Dy+Wio39jNcy8vEhWpvmK7rnfVHOndj1tQ0LbHW/pBkWxxvv5korfoAQlfWXEiy+l
sWHhLxSD6XaEvlvewb7/Hy0a95JnA8CpSMoFQIzKNAK1twODFiA+fYcdLXx2nHPTyw10Qt5ZWPw6
6J+jWak2A33QqpJPUElmUFLCTF2dpjh6Su7q3xliVFSFqRDTO2PWdHp++DQdSCwrynvg4cfUFqcK
aVH8GndmgOdsWZL2EOEwa7aRLRGuZAcu0yQM8pOdd084FyuvD7LUv3b3gWZZGYIO78thOKSBFh8d
H/U+TloP5tQCaVjXJI1yQbpKkNeEZmZ4vFPw8/XDeI/kMr+ttK4g3/ytxhfSntJPf74AIN1NvsGX
5/q0gc5DwpQ13oSNEVsznZPE7wv1BzMAJ1qsqybWUsI+D10Fo8ZxKy466HXyHeqC1Fu2F91regNq
GoYwrnpQly006OwZG8EXj3pgkV2tb2u/RqXVPhIfKWRLH9Hk6q5Qj0crble4f7wRkZrW5zbx/lwq
U43gMUJWinS9HimmmDDvCL3cMdgrLwhDuMP1vt8uGz8PAhCuUljniLi08ce+vBgsuEuTgRf9Zpor
sz/L0hQZm8lfyB+AAelnImOyzxLjAU5J8tWhSk0AapUMy/4EDuyTnjY5r/Ro1MC8q4lBFrYKUALO
zxybFHd47QyAa/rCyzQ2m1k7s8TrG2BFfKb/fYkDd2y20sDOf1T/ZWaU94Vzcs7+X1xvm3u+r3Ys
vJmRfr3CMNr3pS4HLmumIDIE2DnAvQmyhXusmclWS/PxTR+xYfW22DhmaOp8GaSSgQE3g2VrB3iQ
K4CkmLm0aCHxnE7VwaGhm9l0voLajNBy41c8kEhQN0QlmxiXhmp83LAxs7YN8gNC1wwph/+Gmc7I
Yjs4K/7wH7ghJIXxgVRl/88F2FHCAF/tEe2mbqZNyDcNV0hY8FXIPJ+Dw1AT8E7xRQ8HdzhdFchT
X46hizNAHyvIICzqhOWDIRoNbSBzSG3xuWa0fwrWPZD5Z9YDTEcm0wmjo+7tQG/CEQgKAe1GXP9c
Hd8uLczGLt/hWN4re6DdCujULsuG9HGZ1NLgP5Aom3eP+FTdLznMba9z25hblMMiea++LgyAdzZB
d1T8JFVd/JMJaN1TQVNfED4XpxSfY0GP6xw7e/6J47ki4VNpDWCKApI7DklVWvSZ4KS7ndkRej86
EUT6urxch5Ex3ARxqQe5Dyz40i5DJ1HYZPmpVvSlMO72+7S2MVjVtEnbXOWtJU/nhY+NsE8SfWsE
9TVy0Lali/wRRKOMQ5uUEQhwrArwkXaUXXZj3WYbO8SC6eqwt/Z2AV+bA5wi+/4MOHBHviniWlDu
M6mbjfr7XWLBz3h3WIAlhh+v21SPk79A+zGQtpCqBFeWSHVinpd7M2O2mYLUoFkPzD/iWARvbJQW
4G6Ao2MXOrMJdIwiqkG8S+OmIAC4OnHOUsq5fzuXCKkkh7jGr3TpmjmLQYqPCdTvP22KwIB/qQ2n
egF0/VtxF6RXYXOJ3plK3jxT8Ew/PcUxCO+9UAyuLy4htZsKW14bDiI8gkHd1Ks3wll//mp3Ry4Z
pVwZ8eyoRJZgEqdk3DsrCRB7ApXnvIHP1tdeAiv5jhr6TLttp4tk4V7/e8301/4l2f+8SRGRmqvu
MeniBgJ7oUv/QcMfq+LCtyOQxN13q6ZyfliHnn9CMMw8mXuGsuwolAPFm/MlMnQixIWeJOWNauVU
cMJ1QiOceiAS4xqQo9pkRzg6N2j9yC7r2052yKe++6vNiGqcxbESywGrWtQ77DmHJkj9thKtz4xA
lY9noXyswrGbtFB2Wrw2jeJrxE4KKmxEl7m1R8PdXOHQOIFoSkNS6VsqdlCw16Yoy/mWIpvI55MP
EcfenneaW9NI3UoYH2q8mOX8rfuzLuNpSasQP7OIBS83MxZwuMuLkB1+50TUQEWzIT7Em84LSGa7
8vHZ6qFQomhGtrlp/9/l4sVz8rcYkctWOU2RWpHum1H9VvcZmTrxJz2ZY9/7BGkE7EAveqIffLlr
LqIMtg/4blvr7eYDKw4Btory2z3BFCIUiso9HHtyUZCgYhyBYDMZjzbQeEXd2a4tcweJEkMq/EgI
5L4J43h28/B+N6Y33H9A9sJrEYDQliB5DoolgaR/fjM8f7zkD36G+FObZlazESVYoKsfjcY5x67O
o2aCrcvHI0/eQDBBkB6Q7aJqFbP+9A1HFFRhgfF93KCSSh0fIDdmzcWWEKMyE4HLWX2ee1NXe2WA
uFT3IeSQvmrCRy+lnkjFWqAWYrYToBVZJHjIcETvlQGZQ0eIzVUhn/vnYUD6wBTMib8TAwfQ8Ay9
XVdhtOLVAvCNfugSTkSc8G9GK2g3VnaPGUANDS4s5Cxal9XDZ3dahlM+1SgPnrQp6b2gGY3TmAKE
KjI7Isg24JgoPh6B6fj1C3WrsvUj++tpUQtQcfxbUxMNycL01Y4EWoXoi7RaZqeu7+ON
`pragma protect end_protected
