��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��5��+&�'`�|��F�"��dQ?h�6��<k�U�/��䌆�<����W�uV<��?��y�vZc�&�����r�=ȼ��ђ��DC9��Its��<�q�H�?��ٮ��	��Ҋ�v����4�� x�"�@�_�6E�o8#��5��4�f�d��-��C��n�|N��������/
mGz��$|�Ѝ�T�'�qY�!�l�drj���e�%�YE>>%\��E�\]bt/;*�hΚ��wyD2���ځ	��v��	S�\hI�t��l\�:�B
6/]�UXz+��c�<�+<�Y.�'����A�&� 	�=����]w�Rw��=��#�?�:���R�v� �/;vd^�1�B�������,FV���.Nր�+�4,��"��n�V��T�\!+yk-I)�"�����Ir3r���L�U�U'�k�ɂ-B&!��%(�G�H��O���܉�J�
1$���7��Y��x�/vP�T�[.[r7�s��iN��-o���4kG%�$��'�.�s!�m�]رG����)T�*��ĵm�L���"��v���s\��3�^&_��y�k޽5���܍�dm��z�H�	b�M_jl�	�^�I[VR�Id�>f�b)�~�**�� 1��%e ��W�^��Ӥ�MO���9��#SV��
z�i�?�8�["~z t�������,�91����ws[��f��U�ɫ ��F�ІRG־G�;�ge
�@����Ԯ��֙�Np����.Zem���]���^�g�H9e�ğ0G�b#������3����*i�w�g�t�,82t�oL*��s%�1���L�RN����77��<�o���;)�5O�&� U��t��-D�����uTݶy���,l��%��M��>Ɛ�kn����y�57��Fo(ʀQ���B�f�zk�	���E���'�Y�K�+�o0�$�����i�Z�4�3A��V��7��p�A�Om���g��`��Y�^B|�6a+�13E�l ���I`��!�0Ɋ/��7j�[��υ-��>�����o�%��[��|��D8i�,��V�WJjY�xUf`H�}%I�ЬNU��ȉ�^�\"`CwP�M����y�����i������n蠟j�%-U�m��$3J<�Է���b��E?�����i	O��1��P��l/F��ߨ�!��*��S[�6&�3�������� IM,$��Rzϑ�i9�F��|7�
��.�e�v�m-oa�e<Hĕ��_���׿p��|H�6z�(q�R���R�-����פM�����0%�����,:ZZŅ�*��x[M��ˁ!3Y����-=w�d�F6]��u� �t��0He�$7��߼C`&��p�7��:�Y����H���|��<�����gޡ3�|��LZ�f�"<��{Œ�}l^>���a��+�6��x���z�W�2�2��`�T`K)�G�\8|�iq5�+�-�r�y��XӜض3��O~��$�N/Ӈ����0����n�u1�x�M���`�7�����ȟþ^5����j���aC�g'�z<�5�R�h2�OY?��㶵߀��Aa��񊳊��m����������ye���Ɋ���^�5@�P6��{���V;����4��&xem�]M�Z���w^�oy䚠m�� ���+?��漢�f�dU�����u���GU|����4�*6�: 6�FRE�<n��C_������~���/���2|����M��%��^��Kk��� �d]�?��1�Qe�� �1/�!ӎ�=�,�	,�յ$LA^�[�ǻy���g���t��|��?M챽u�
]��'���6ܾt���b����@�n^�ǂ|<����<�����Ɍ�o�S��b���@{���jU_eR�G����X�Nf���Mtfd�r3�ڔ
0�G
�;Ca��}�N&�Z�h������Lh}X|ڡ���u�Gk2T�������-gQz%G��eusU(�Gh�p5 ���JM��	�WM�\�QK�Oke��&X_��K�r��.�ۢ��ʠ�	��(�)��?��c���B_&��=�	�l@�蟎�� �I�`���z_in�A��$��e~I�	#l��nk�~��nGis�Ao����?�U��5s���fMz�t���r�A�}��6f����N@��b�h�����b����=��ýB_e�YN��)��Z��x:F�=�~�� 9nP�li^��uJ�����ص!�җ��e����lS�\=Q��v����أ�=B&� 3"�ϫ�����)�Y惈���q�iF�ƍ��.���]ّ�ى���k�7�c	R�,���OJ_��4_��s3fض��#�繭�D �ڡ1��D?N�K`�jc#.�J�1<��q��ք��L� �-~�R.�͌%2/)8!
s��P>��
/��L'[J�E�{-���+kmӌ�k՘��ִ����#�1ݏ��;I4>7թsHD�Lԝ��gL��K2+�;3����Y3�BpK�0J>�&}X��ճ��p,k?伄'E��y4,o�|��`����ӗtǥ6��V8�<�ŴJ-H{�
TF�'�`j�1��}g~j&>��\�s�D�wG�Ʋ�D߸�Ip/S�<����y�vn���2�휒����ƶH����lz'����:qgܴ�)�MЄ�tlmg�ݠ2jU'��ġ'NbV)�1|�*y
tJ
��L��}[ӑ�w ���Ħ!~3�;�ꡞ6���P5���,8hSRl!W"���Nh�?Ũ������_�Ǳr�S(����u�d-�Of�6�|��:�8+)����tS�Ѩ�~�b��g0l�0i�nefuA��k��C�L�f4T��7�<_ji(i!��M�D�����i{�1��vK�S�;��3U0|^��s�a�*v�ь5�qs���f�=Wt����m!��0-���#�䗳�U�����QUޠ@��F�1�F����p�U�?�w�t�poOEp;x�Ë�����^�yս�f�;�z�^J�5�Vƹ���6�E����E��Ʊ7�>b ^���!�*ō���S��IH�B}]>���p��'�A�J�u��47�K�<�����;�~�=�vKЮ#Q���y?����c]���y��qv��=���+O�����02:︋`��g�������hR���Kس��v��B`^uSO1C�ۼh�,@4� �RĘ���,@����`��E)&�h�4���]�1�I�=?L�d�����73���Kn�Ar����E"b�>��EG3���B�5Ol�����B�/PD<Pv$[�}����M���x]�����\���" \�M�ֆ���*G-S�I'���I�v�3?��$�@b�O��)��	����_&�BA� ۬��vG�~=�C1�nDi]��|%Mҍk�Il�tn1v1��HԷ�����a����z�����$�hf�SCU�-K]Qn���<�8� ���y}�!��{���n�~���t\�������poV-NE=:�����uIX�?����z���������Jc�q�ɀ�&�p�2%.!D6��*i�#�y��q$��y���oti�Bѽ�����au��ۿ�&� 8X׳���i��U�>d����d~�h���V)�X��p�LEi��7�K1��e�<��(N�]AOU�1�K������K�@?���0��gN�#�կr�qL�3�e�� 2��4&��a>���ɓ�GX����,T�U��C]*5jS�6>�E��<#���U��ă�jn�{�u\cx��V���/���3����M����^^Nə�G��w�m�3�GǕ�!�:��º+�w�R���ϐ�Me��>�1.��N��=�a���|�T�9�SE�������	�+m���T|����=K��"	��<�6�{Ḙ|��>4u��V��{�.ąT��)áվ�L衽,E-1���(ᚲ���+MM���pТך��T�b���^|�T s�k>U�d%iV�#H���z�f�V�#�6�H+���n�艶�$�,���f#]�JH��(x�TOv�yT*��Ə�gm4��!�y����ޚBL��iz�w=�<�at��u/P_Y{yy�������X���O���~�F��þQ�Wͫ���i-Յu�����F�=ڐ�t���͹�j�
����7�⡋�]/>���@*8u��â�U��Z��$bNf�k= }_Dk/7*<��*5.�(�~��o�e��ꄦ�Ҭ�7uAv�/��T�p33�S�6��[N���f�22W��EZ8�b���ѓ�VV��t�VNA弁����ՠ��ڹ�ۓw [���/��a��4����uKC�փ�2�@�� �t�}�W�����>}[���d�L�9���t�9�?��T���PQ�x�rk
�"?����j��̑��K�����4cW��8��.�F��gD�&,�]�����/�e�,�XdrL���6)���r�,�wY��$W���.Vo�B������Kwc��"���}kn��o��q���9�3��v�gM��4�����i��a�E��o����W�;��
��(�1X�
�p�@0.ap���.�(e}�9�ٳŖ�9p_ɯ{���8�c�Ϡ}l+@���:��(�/��Ve����0�(������I��[��_�w�J�#&9�Z+�srJE�\�5�?Q^j0���Xx8�7_���o����T[C~�mD����3�y�:�|�9@"��D�\Tʕ��,�`�`*����T2����K@9HF�KVB�C���8�,�;��