// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
UP8pWD8vxXFIOQubecOquvCRp3lWpiCpKbjfSS3Ae8Em++OovXCRLsjJqsCi/jJVdQ7e8yRRsNer
DbT5dATP4wWsZF6S0sPWuMp6x8uY3gYLcCnxTNzB55yhLlBGRkp/bJD5GrrBrKnQ12uxQ3BZT3Gm
SbATlxUmivRPc29pagndKECWOtAJGvFIHP5ckwno2E5EV8EfmN9iOJyeb/fMiUhP33x/t2jwUo7z
yN60w0YkLVmPp3LaHspC0mSpa5JYUcsdL1PNivRC3oKF8TJ9MHYuatmNyBqZAkWIFYRVy+AAeU1c
h74ctQKqYaOdtQdWFLPYEy1GDJyXRb+iBQjbLA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 64880)
BqCbWXEwC2El7TekiMLTYeQiTYglDnEz6SkZkXBCtnL/xY38am1WSL6rIgOSYfDgAMELQI41zgyJ
YjKzvKJpGqBFtvBAsT798r0mw8SKuAJvSUaOoofcRcyCPghwOVLks2U1baHiv05bN6KEj+5zrbjG
FcUW8/EBI89leJ51YmRLf0RNMiVNtELNl9D3NMXtpgaF2Km9GFi7rpdZVjDD4FmbrBo1C9h9ahyH
qU/dpoHszFZHIoT3zXsFwwIO794O6iR6gqkf06sAeEuH2OYn7nM5wCIS0bMMeMh2NH7l8v6A1ks0
jJi10z96SP1Qt8lpcp0d8YVVWmQDC5GJWm/om2qEojRTUROtRKfWap8WZq+Zz6QQMMaXzcnMTMlw
r5BZ74YBO8o2RRuzBdhAvT6rQ7V/dN5T4yXlrocQFb8APQXFSNvobrH2Y5+snRGiqhrex+IqO/pO
r1vJKaidpLraVvqplxTNdzhr+AwL38NVYYNq992Y+T9BMYuFQjieKXUWsykpOeF1ddCBGH9QM/+0
+IrfBi3bQLpvxzMH0VhoylV08WJfjc0hZ2tWcJwY7jMFxZevXBN0LFMVjfSE//2oVRxp1QQI4uCy
KHMsyg5B73GadPOMSfZ0lq8tFKbiNYexr2nYhqoQq+L4mOEl9UybCrujqb4vNstpnScNPrJ+gLnE
IESjp5/eyPACFoZ7q/jLAi2x305DC8MX3kFzyTt2uChVdnvplKmxVc/L3a0bgIlJfjw9EO3a5UEv
oOHNagReFdr1W33MJA7LnZaJVHZvWJW6AOqvWhtJB2TMG4MWhUiXbfg1BV5e/NEIqrVgR3XZIPxq
bJbt3NNCZ4cJarCXwQOvo4n1ZhSz8OtChUvzO3PLw7UstLxTZ6mrDwmHW530Urrx+9PVpsN7Gpot
V84lyiBB8kVWo09KTE4n4xEI5Z2VTxl5ZNDd5SWNmdxkXw/+Zev1RrUIZ/YRVgNHulbTBxc9JzxG
JfkIhAdj8CRH4B6b4Wk8PSFBZJFTsJaHH1U7LWQM/XqnFcWBr2S//UVMEzifYqjpfA12watbJldz
8bZi0AuNVgqYVaiFAR0PH21tjJhs7lr1/jCaLHmaloXGpM8vYkPzmvKoRkGvo1R8eAHz4vyiCaF+
KYVzOfQ82hTv8/AwA/VNsF/99FG90exdatFOo+0MkYCz8orNPZmA9S8cwgRVQcqk+Gq5hdLRkmAb
uroC0XDEoZeVMr2qrY1rj2uLvUOPgQnN0/DRKShyUKB8WCIxFXYMdQ3EOajOprRBJS/Vv9nha/mi
QA41FlTwFwuebay1U6LUjtgTlGx3oDfMZhKzphh++UroN6j8ObfDZLT13hc7dZW4oHRSb2Qeng2Y
zrBF4K2t4ADlYkYJ06pyP0nqFK/+7uta2ETW2wnSGJjYcz9LG33d/nWOMlETTP96ZPd4Oqcnp8Id
yN5DpP9yEgCYqt0S9krHOyUPBuXgIeTQPG9Sg/O9nN4zD3u70xrypxMK+rUJm5MO/7Of/4MhUO0H
apxtsay4i8QCFNj96ED0cGIE2mEMywpCZPB0jENSHlJQtGMjXlY13SDEQ+6L9c0pN2wh9dfL+blr
RhvsBGK9PtQHHOC4ZckjJ9lZMhN4c3Q6K/RiwxiqfFnUCF0DDlDR9mLWW8oCZ+Xck4zWwyeXdUD8
eNfn9ZDhxafXu1bA6WyNre+J2QkhltvBt/dOoXTKzjiGurtIZgkmJ2JOvBGkdz4a9x4oVJUdN8tk
EwvQuskoCNRjlyH4neKYt4FTZrP68NbUITInQGJ3MGq4532UPFt8pWVkO9cOvn7BvmYG95HOaOte
V1sb+ZtmthpX90o85jfdGTELf87FuPu1H156uMdfLpvlRA2AsXidstoNiMjXs3una6SJouxmmZ8y
iisgVg2gUrLgv6rHKmH6WVrO6rAndgrG5dUTRedCMZj5xATnEX6h1p4a3H0FzxGzRZrctonPvGNy
ygng19tbEAEo8w2oC9M3AoKs/BrN2D0PPMT7tk+BtQltG4RrGSmdy50hdX1WcqSaRN5Aa7CtrHk3
lSOO+bEL3MgsS24pnPCzjXfLQ8Q06y77JiXLFsbtHBOR+15M0gjMl8+i0j7YcAhXhKo8REo/o3MI
m6jGiq93bXhPg9B35Vc1EC+S4x2IebQ/pFdm8C3QiFepsJrN84tXtHiWsVAaKsLrT8PuvnCuFMbA
l2V+gZ5885WjtbyvZzQtc0QEZMETk1+fiQ4AAgmufEY0eUI5020c0866MLZ+YDlJrtf1fXxqvQwX
1kMHtCYgnXrHoiBScs7V9r6uS5mOr5GMoMdn+/LUyak4ZdJgG6kKhcBweFI3dIxDzay1edGlzfCx
d7jUgs/5l2cFJnO59vcBIW7Bk+hJpN1nlnQr6zYEO+OzRXcJkWweP9OMOPbYnEtMRhTc7P3nQAgC
OGksoUJ6PD0t8DrwDd0EDmClZanJX6cUsBO+8LVA1yZgDSpOxhWZDbg8KgCLc//8w+PDl2ShtMB0
78ZG3mWUNYuewTP94+ZhA5d7pFIrisPGbWQP5JtXQO1hKcOOhs1hgQYxCdU9DuRaAQSaFjQBOgY2
VeZg3vQhVTIOF+L4bmsuvNcmDa2A7inSGfGo7YkHnzi+j4U6Vz6zSDFcwpFQQ1Z0/78k0CZsxQkD
UjIEIfMtCWF8gBc9I8V+jciKJ0BFwmCwkwwFIks4C0uh77mFmT0VDRKblsDAKGx5kdhjQvx9XYBs
R4Hq1elK4Gctmzp1E5QkvlWJ5AodGZlHo60Rk2hRR44RTIbKaNiDN8I2WIZ+hA1HgSxSj+tyzwn5
ubll6Dv8dYj+fpQnE/ZuBuj+eDvMw4yffm0EKFNQUN0/wU/AwyjvTARXqm3mf9FzvtIxxxNCeF9q
1DaU5o2to+VRWB8KSFz+kEHHUFypQYHIVWspO+6NK4V7FBJ/jkk2GBqo2KY5A28gJr5ZMm28q67a
EQom1pMnuWIQvJVIJSKZDNAKpge0/aplpOXE0vBEZKEXBrqBvcjxukAnB3DfjJeqCrPxOYCxYcif
QVqJCkRX0OJmN1AZAVUxGqLj+2BiD1bswTtCniXj8k9YWe5PVpUgjNAPXrhm9LlO8/59Mnvl4c5n
KfpKdrYcmy4WipZO+dIvbrBRBURj/ILEPZDgcvWPubcxjaRFdFwCrgd0LZtCgWmN2L3VX/xECLca
s0fAD+jYzT6Lj77kXDY/+vDmvqJpnzSfShq/vdBzYIAu4q6sfRCyfx3sxHYMEINsN+e15Fhy5tOC
vyrF6F11aIbavQZf3JMxzc0eP9R5XrCLM+XYWBkWd5eh+rnBp8i7RPKb85W8iD+fYWNkrDAfxu5s
inKOC9aBktpFPz0cp3DGxL0lwhY+PyZjE8nsequjgftvSXp7x/wmF2Ufg0gnOJ7onM96GbgHk5QH
a0LUZpr2o3c5sYx3Tt7y5523jl0HHLJ7Aa0UfsK+VFI/rxG1AacSCVAaODZdNXk/CAjqCpPgF60h
L+Q4A8FhKOBB223SaS32YzAbR/1WgsEiU6J93sn+T/sQ9YTDi77rNFFMixccx4JmiMvfcIfHZ5ys
7GaD/mNysjWx0V/nFYEt4yTMA+ua0eZsvPRFvNTjkygSkD1s5ebpJF4u3zj0ZvKZe54fux9S9hJK
rujtXVN2LOlvcy7HMWIfhFP4lPKVU7IS5GOBauTQ+JDGvrUuGcbY9FrBXi3tRYVJIa0Z6/3HhnVJ
9JUrqrJWYuNoMcmXjiZO6ffPvOrqRETaGIOQXkgs0dYnyUceI9zTLCE+BbzDhIzkdzxFXNAdJVAR
Nn6zyKNC1ctd0GmkkP6VSAPVYsvEQ8W1EH5SXV9G4IRPKM08JhPs1rY9TZj5XcCTu6WaE4CwqnZf
w25xeWucBKND4dfDzwhnA0ZwwzUCoWpbnX1WQjPWRAiuORQB8mjqKpc3K62kGPjViJsiKP5VKZVn
EErMtNWbFG7+bAeme21HR2fpanLGoGzG/bZQfMhTQ/6zVAX9H+EsZonwmMYpok67e1v2+W+b5RU+
7bn33+1cUi7lw/im1qOoRzGt7oY7s5XTJPnQrRpsyGUbT0S35SPxApyn5cuWYGdGG+Mb9HyP04sK
H+VmLC0CkKU7oXt0NdjJlwCffrSCCCSKusM3+RKQui3c+dnPsdiEZTEcX938I2cRbkLYGfCHztRc
r8y/5zoStzLjitL0bBPeggzn/ocviR/P1RO26yQlrq90sktu2RVnM219ULNuEE5DAhlqZu82suwb
39UdgYPIFjZSAWAiRQOz+nEzknFqPGMJ3rwWWBkNkga8wKuzhZmkRA+ry9Zsm/mTd/VhzJT/qZH7
2+er7sVtlS2vzKusLprfXfbygxhwLzQmM1VzI/MQ8xcJburtWXoMjSmzZHJ1ikgrVa8t234UwnWN
jeLAXfIpGnHyYRpGTLTbCSOGEmoVjTRtUZduRQYbjz17T0JxJ1YavnULPtS44mJ94QPivMNzatK+
Xdn+8sOX1Ida5PUZr7Iyr/+06rZcN1h8wwnm+s7vUBwXSYL12l6avD6jCbmGwfwDkvEGnYm9GxqK
iCXJPfwbRhwW7E8VtdSWm1hlUG+wZWuefcUNsnUAxuvA55j9HKXhX9/kpmjdk3bOwBFTPT3qCQe0
QjIK98gGg4EUFjbJBxmZs8RMAAfKI1+Xw/4V1QwPQ3PReKPRIBtj1+kIS0V65+npMc/1LWBNpHKi
De9Q7Qn/RCwwUeIqZx3Em8bLlgwivJ7/6OQ6GFhGBeO21YKV7YT7t8lHfP5ZjED/qNJp1tJAPOYP
qJz81pWwqq3rkrdCDwzyP1syEh+Dnt06HCPz0drZpswhraCD4wDTJS6+X5vS9U+a2y+ewQ3QUf+L
NUu/+vq7iKfNUppmj420aJf6sI6b8pnFQRDItuvm8VZSV+QxS6ddhivQAc0y+SLZJKAQMSvQqSRD
HIYx0Ue2QULOyhSuco1JNdr1pc9OseoKrh/RpZHa9AWg2jtBIgjC2pey7FTWy6wtYriFeeV6s+LH
ULCVUcW5CWLazSVQoNcBwO969A6JFjjNd3NBkqJi+yebqq0TAnfie1JDYdcgxNtpvfMdsvR2hhub
2I0qqS1tNukOH062xxODG5t6XvItjJmgEeVZbq/8Y4oBsADv74YfciyhvdXriShOTrcD3LDu4miy
3ndttWVhL5s7I5gjBYuJ22Is8aflnWwoiN9adB+bQMYuF2pWGtnn7s3/yXMveokR7/ngWBRfB1Iu
7miBEsS3tIq1dm5tltEuLMtdz/n0t4OKPNzSnQrsNUIlB0ERcaUJwQfLKxmvaMuC9mbXRMWijfyc
i1CwamVrxbh1PkIVOEsX9BhCAOJO/fA9EjCeE6C5tqMane/mI8oFg20Elg1QiPdvj/I1udRcbjYZ
I0o6jUudYI84y8BTCkHzgFHVpItj3JbM/4YMVkXJreH0SjdUWnjLK+IN5ZYKu38KjbxHD9ZSi9u2
lq/zUtgywELEcNd6JYszWsqnH9eNCpYVgz0XoVG1RCc6e/7WyworltnJQGtNOSeW6VRLbbuH4cdd
Wto49LmBrbHozr/N04Dl6LdSW/W5fQ3F4xyKXPmcNFoVN/xSKiFX8PblCMtcJ9xwJ9EI2EhvGOvM
l4ILpCnApvPoTe2LVXR0hT9RSS9jFsiqs1hyWn5Ivq0upZN5eZhCPoBd9+g2/cN0uhrqsBUgnsuB
i0xPQeXNJgjvtc88+jtnowM8kV8+aJu6NWCL1/MYH7oxwQfV/wUwR8Vi4mb5W1a0xmY39SmUQA7x
XKUY9YNVKK7aMAnu2o5Q7r8jnBKjKqa6nO33/e2JtDq+IN+h3Oq7/M0B2qPBR9MNay2KLyJr7ldZ
+KENofcRx2Gd9zxNJeceHpuGUj5poC4BZGQB1vQ7jp+ojz2HlyDV2LXDIRcPLQVfJIxpFRTulQ28
0V9hBdqoNDcE8J1MB5Xbo4hPQVMtbOqHVS6aokI9hyuFIZHbbkCXN1eJqEhJmrgkrw3bo0uA5cgV
n/dBquNFD3dwHLUmCHXmdM4m9n/G91Kwi8EYrmd3mek7LY7z/pTSAju03hljWWqfxs0KLJZs67EG
YxuhFD3oZtKDGJUxYhf/8QU0MTmfcWZffFtFLZ7h9LsH5PopeHqirUxWbq8TC8ySCmJScYCdz1rt
ta7FWqlNkMW4XMs9lvCcTuNxf606iFYpKRddUreY6oshG7bdlXP3iF383I7+4cv8wpI8DI04f8VX
8tWCTpg5C6WKOm5kNock3ptpDkXXsXJJKhLn4eRiFLQWBktmB7bacdCugwDe57ynwbt0bCwkGVyQ
wuYrtz18AJPhXgxR3ukAEen6AerSM3nKGTNMjqWeEwqXWOVJsLJero61ijeHEqVGpPfBhkyQY9n6
x6HM5dv0Hrnvan8Suqb1WtmXuOdUqNhbFdZtjmgMHS601XX2wI/2CBa4JpheTxjGyQga12Xq54g9
mwrc6msKQ9LLsEc7Kz8zKzgy2pqaVlMtVI39mrdsNvdilGkdL7GwUqWr+c9NlZn/DGP+eIlv6opY
s/xYLHFUNzhFwT7PvHTaZaA+sJPd4GQ6lRXCmo7GmoC0lBLIyz4uCkucDz/xYaf9t8jblLvWaHf/
7aV0o9jBhlQzZUbMvorzf3bfhpfcdeH9KbZcvqDqpnNPnU+s5/LURv+zyI+OAAMyCoe7d5SPvknV
55a0UqmJVJRSovy/Eyd4y5S6je/ifzXp85KhJtc8qAmCf31EATxwfSOZMK21vc0g8JDqk52qKDdc
CPOE1BiGqG7CLm5kdJjwvKuI1Hcc4+U4Yxb7nC02YQ5EkLcZPtj1RjMgHuNJPj81hLsb9xyjLHR4
fJfy01GOZLFzSNz6qk4Wkx6OlcsfZYYAdJas9DGNnTZjGqh/lg0H+XA/zq/tf2uHq/zjJm4xdvSi
B7cIf0zduy1kJdWqQ4s0V8YwDsMwqYbMcUfWKa6/IPjoOKIE46gjPWXDgN+tnEL4QBpS+olss25F
F+/vNsfC40W+jolxCZzx2DB0xZIjWUwhhahedjAYrvJ4dzccw9ym9Wl5DUjEkzdXUkfRVYg41QV1
OXI7t4nfCkX4I/yH2Nh8N8tVU2FXQ2iuHKrci73dXE1zszlvIUfXcwNnFuaUGb+VrrGBXfl/VK+C
vb16USQvF8aIuqmR4cLXGETVnCeMTqFA7UakiOzBv/FOIeuOWnn3wuHtceBS8QSlVcKFnzB6kJDF
qF8ciiH8YoAjLyd6IzHDz6jsXOAAgm6ogy8MeoNHTq/lPy47n7zX4gMraKCDIj/ZQGMl8kJ3UGtI
4luQWD8nj9n2kANIlVewMtRIK3svecrO81iLSxe2KkDYX9QfvkHC8wjW5wof/GDpm5NInJc5WhPl
4nN+BS3sdFN/UKMIeGCgOxbI3uI1DsR509mKyVpkGaitOrpZH92CXDEuYWMElwG0v9+9uetuDT4U
50dLPFdp9sCGXo9kqrSHcNvbaA9l8kkAijp59yd6MG3J3YkpWeMgsSgXYAbO1IwhfJ4XC6rLXANw
MJ/BeaS+Ozbhb1emkdw/QMYb8XFJ4or7eORTVHCEvoAJMfHiILAhNlhSZOGVJRnl4vgIPJ3KvjTZ
TWt5c0A0AGuq3f28gvsaVlJbmOYQB511riCqfFejCFlPuT2yVyfXMeBUUpEjWci7UM9M9EmzF8nq
GmFX4wzMZhyeCbhjWCW7VgmkOFcF+P7y+0qT8uFsjLLAR5Q4qOb3oBflxuqFONhKir1uqz4l/Ykn
r4+2UhKc5Fq9zY6ZZcM0kxiL4TK0TRiYldGgrfhc9oMIkt9CYa4cZMjQnP/D3fcphEYkeGOH3rO6
P0n0vMC3LkoPKh2vkUr/fvx3/AqmSybGaPN0ofyV+jMj0kbVfL4VxMzIT4gDRTCtgoZ8Gvn6Lv6o
3qUiJSEMWUS3KIBGze1PFP45Es3FosWGeHYXyhmDyx4CR58oC5J6Oiffd68f5WJ42IbrYZ/ib/VA
hKt9tfbublJWezs8MzDLkUIHMTuZD4LNG3c+b/EaeAuKLzRKbpy04C7/klTxmCJuZ5MmAlJgEofa
8jJmPrVZUgffiA7kl60aWIFbPWh+snMFuMVSjULkvQF4qds6/HxHfK5gGk0/JF+lPQjQzkch2tuI
M7oE43YaYPsbtcD+8I08WFXa2J5jJZ4aiRUAmLqdYRLH0uq6Rp3s44C6GuP+7XvgA/EC05w2WUMW
YKX3VoyXg5zbTwx1JYK/408ZYhQ1dImivtlXe9CN+64V6Mmkw0q/dv+nNuQh0xp1sFPIroI+u6ng
0FdCD+jhQWOd9KOkyZ9RGnrsjTeGq6At6mW+vb91OErML07WrZeZeCZsj3nZ8xvxoXC4vb/W2bo9
EKFZPPFE1UlPUcCBVq1nB7//DRsPy+8t3GmWCksE3Lsb4jM2L7Q40USkIOgvrMdzBqp/y0pZG0PF
97KaCGsgf/8Bc/3pTwKUUqPL+TYeUbX5sBc2zaxN0OU2Z8HSwGRpXKo1rbo27OzN293HUS6oP9tL
1xq0azKZ/0FR64GhgGW3alkOTDlNT67tX31Z0Ym7wpQQVIM06yOwpqJL1tgf4nUeuwPBOO4NnGex
LeQZwsY3VXJivrb5werdaXo3xAObg+GAMUEmkywtHPRWF5zHxjN78DOQmy6wyB2oEISM4LNVloVV
LHfGRyUS7KeR13UAGSquotq3qFpyr7MNph0wveqFsWK7NkEVNRCbHwv/jKXZQlYshzKiHjQ3bY5L
rUdE/aDu/17A1YDsdfbNMq2T9alx/gCroAhR96WVYJmO9COctanILA2jF3Ul7e7Cc6oKHtI6i87z
62cgAxKUJzeufg+SDUzkBkXKJ8dm4HE4BKOwxaqpdHd912Z4POYS8wIPLlgLmnVqB6DjtjZni0e0
qOdwt0Q78A1AblXA01mceJkoHayMkc/3hlD0J2My5dqXqyKBCEBWHwrjBgBUpv+FA2/PeqzZk7NX
ZjtPXvyjapnQZ4X2ziYUEF5WvJt5RyqhY72DCRNSCKJ+nST6yRDTtlehKfbzCjPa8e+KZru6Bqcp
b0DZsmvOKS/nqAZuNf3H6YKSQuBVxXorWMZzzSF8xe3gaQKPzbLSvVt9c0FAPBxWH9sTrFmtl6DS
nFxeFRcbOTrpnEy4A5NwnA9PI9qSDe9SH6XjQELKXuoTvjaS+xqIgEk7SKxtvyDYp9N+9XMifFk4
4ZZcEylqvGy294jlS+n910MAS9HEiNSjE1fYijgLl08V2I6P563gEEWmZCgL8haj2deThI6QgHvH
tpZYjEiOk81TEeT+vsK/sZ9Fy5CjNjk8ldv0Eq5K5wmv2rS6ShjCn931IEum5rAJ0d1h82W6zoxc
DY3k6WsFYfS6epvleIoE7Awi6Cm0cAKhGQovGHYWnWUycLVDtm9mCfASXblMfawj6jMqqE5e0Fdo
jSjrysqArc2eDU8Ty977UGeZcoVQih0LCIUu0LwAkECHBPFDGhAP/VSF3dS5ubCrz01AYoQGP35c
ed3mAgwQSNYf64hUrxZ6zfSrU1YRdmlKofKgeMKslJUbvw9NC2LuL3jmBmPhYwZ6evSzrKwfDy3v
PlP7t3cOu2JAHH5oR4UbvRehYNihN5ZQxuDtGEhs4VvdL6180/oQbXtycXiyDu2ZF2WxkuSlismy
SaQ6XsB3UUFa2WikJwxscrRJnXKdBJIUudSKF9f+ry2jzbdPdX9DhU29SBFrjU92BfN4MNzOBYtS
o04lc0Lwfdd0ycTdYiJKN0FXOn+lFL8IPPXxuBnZRfCTPFLME0ZNLVzg0bPR2O1xhR2NItvYWego
7nzwi6kqLszvqo0lODeyz308MkVTS1bI9fEDkmUrWNlYsnZn49wuFqlS3dz33DiFNfNLmd4vlJEz
74mX3Cw+nVttgicrDPAYVIs/FcicBy6RnXV76BkgOE6KCaeeKZ0uPjxyIgSRdrMQ9XWuuMHvU0Kk
2uIAtY3DaU+fgrWKMttqeXC/6e6pfX52w7iAnhkdbS2mnKeRtjWcfG1qiL2Fil9GorA13shSThdV
qSJGhOz+VUnduotPI119ONNLc9U1eczPJDelCOXeLS0wTco1icJG7h/97to42zyQ/19uYtY0KwBD
hiTXBZE6j53Gjuq4rhDLBoZFUcsKn8VdZUi9eP9PcGNsN36zEKol6Jg7+shLKcjak/eCo/9YWZNi
iQRqjJ2KZrzFImekKL2+JONnVMOKU8C1pWmhqwNMsUfcZ1bS7pa1saiZYgl2jP6JSl7VSkMfAuQg
SKuvx5vXKdEPZ/ifgMnOs9YmliJQclCXkyeWMeAitlLgGevQwvU93/3rsWTKFD29+ze0M0XDAc75
QiRjtca36t8hqk3mG4ukDyRHtKmAIZwIHyGQRcUQAONf6mV6qcklfck9Z3uiqhpbHKMqyH/G36Mu
yGITPowP2UdwcMbOHnlEXhKGldkHGUMOgrbXpPS6ySFRsQpPOaCj0FnPZeXgSV5/wEzmqxSIPGiK
1vJgXG4TmiXgVINPYTywsURtN2RVRBv5KkNM22OKzbACU5UNQcfFexTRw7ACZjuTHbPiWlMlOdJ+
P/sWpL+QUmawqsYeb2lTwKN89xTB990DY1q56GuWdHJw/7ALD9T/frFrL5UVSVbDIWP6T8JVP+VQ
5ZJ9H2H1s2yJrG71gV8WUAhHaOlKEzTEwbY/zv04cH+rXAGSS/e5jAisOaUeBLdiNVEyDAOUKH9K
rVk6XS9B2UoJoa06UjysNo0jzWoFvVkshSSxTjOFg79V8MJWmTUFEIFcaZhiatDflyEZSn9mQHXn
vV4VoJzlagOcmcUIrrJLL6Xlh5Mw5LW7G8rHjBhDuRq0jZqJ5jRMKSIV0JTbBLHdKf/hdvFHk2Mi
avTAV1A+tcOIfjzDngZV8GX16BaXZarLTXYT7eiLeNz3JLqiCfihN4kxyU2DjZST2mIU7PiO/e68
TqJFcfyjjRASPwVd+BuruIQkLgqEFNe2Z1+fD7SmCDjv4VFXYf2uTQvTnqMW2IAHryK2oGocyiWn
oTyBzTER40U8Glr/iS/mgHCQJ4z0rsma2bs72TeGuLFMFC0SHVDp24ktg7HuMLT/PUPXRKCHkHal
655jysa8laAjG7nQfEylu4cJ3A8xx7oENAxetZVL35aWHctXS/veTGJtcU5EaV08SqUlDdf0txXo
Wz3oCS+5t5wcDmwyAUeJ9CmaAI8tPpJXM2me4uaUgun8Jn5Xod0Qvs4PVAXeqXWVLPQ4dKDrQufe
Qe32vA0bHe2efdiOoo2+yqms13TneSmi6JOoA19NMwfHQo3BAwn9domJDYPo/hDghv+ngIFONBAI
btQpRUH/zivnzUbI1dZymsHBbQJpyIIO0ZHRJMqfqZGm1M7oidXHDdXluj5RRMH00N6lQk3L+yxJ
1Wxqjv4xGCdzzaOSpLUlNNnKcssKqTIyerssDE9FeNdE9OrFuolhfyj8ol6I7QZe015KgDEzJPxc
1EJYYKCimcjqgUyJ4YRtvvns7jSLWgJ88PCmHJziBs2NeysL8vx2Fz+/pOEwgUDTIf5vKdgW4EZv
6Nv0W7cLlFWM+wRRVwXf0zgaE5v76h7taxe/Ic1Q1EDzWcuRJtDkSvKChiiL0+arkHuwLe/XhK2A
QA6s5oVO8iwe/NUbVY2m3k5lSt7ZgTs/lmOmLpM5N0qzWkZZFrlq1IlYjsfodEk1N/XWGcq0hi82
yBkQV1RZe85jHky84M1/4UjwTDlTuTtSexmxjZo0Kzgddrt0vuRIErOi48HBmEWBpfDhw6E3sMWq
CBfzI6G3/nMbPVu8vHizk4iRk0oZppGuOoU4H4TYJcaYm4r9+usdqa4b1hQVo55/hQeVDfaR8oIt
lQBkq9tnctjIIbOPKRlEC34N0Wp/jGe2N0KaFUmJ5EvqdJIbnmP6dXo+vi4Pj+B4iUwxMl9n10kn
YLHZPGhCNWMWi0jroAaEIi8VI7g1YmTt3XXdhOEjM9EBh1+MKerzLx2koWg/5a+9/FrAbb4JNwIx
LrLfIFhCjXiXHTVaEKClhugq48x5kLT5wiIy5NjUFy5iKFLcPadQxRnkkJApxkGsJb8h3JA8BNCu
/Yx+hvP9XesOAnJ1yYYFJFBVLiBRnxpgvGvYTCCkkQSP7ZYo9JuxczReLYSWDtnkbgvGiPSS5X3D
xUHAnh6FCSV1gvhaD/OPgAzlo4+ZQ+3JPYq/A5867YBCq4yL7++OmQTe5f68rpQpBAHWEQOoNXu6
xk3Auwl5cNuOt7YwjH2EyH7FRhDiyw6BJs+hkcBk8/WlXwVuk2N3Nudf0PXoGUr6Kni80zP/Aemc
iu1NpL4emkkDpL3uVxojbaLF3NdWT7y9s9BHLb7d+p4LkoeVmRBsmtlYKinVgGHiQrXjqv87FeMl
tteFZp3lpkoUcToNBZAbqm763QRoMoZpYW+youBamviROAhW6EaToT+q4rwcL4CSUzNzK8J3h358
5macW//uVVFtL/1GfaphJW0y3euIBL4LBiSNCC6TWe3x/sgd1gwZFrhxUBC25FHBoDg98i8ro8oP
zuPhoT84NZ9xjBCwBqoGtD51uPi5zV2ju/ZbMRLxm9MewhG0hz8jx4awRhFwllISrdXWPu7mOQoM
3twj37mJZ0sH+BBIVFJwNzZFFCumhQX05qXb0CCnFBvRk1ZcVBRC6fnpTuemSmiWrVAk2K4OUuWt
S41BEoD9whBqaWmMhdd58BKT4n+9VqladC9wfNExq/4lM9BkqJZGNWS6Th7V3PQkDj7FXJ24FS3a
IRxnL6fiIA1PKY8W3ojrdydZdxsODY2Y9pLWZb/Fhf0Rf4u6kyWoT4+RHA/WNE7xqIVdyOFE63F8
RHeoBn1fdVv2AfpA02KD5zoJ8u/MkHtvhexWjSgJtFG2+RJCq/r1W9g9daGBJKGgRoNPxJgEWON4
ek4s7SEqTFsFaLuJ+JJCjqorC5nOnB+JG17XOfDsCZCIe6z3URJBYtNkYiS8oOlVnKtUCoy6arvI
9KZPCj0vKpGA+VJ6Bu14cRFygWSGv96pf2q3J6BBiY6q7G8LMrsU9Nuexi8zZ8iUwhS1T90mzwi3
bsJF2tsEk308grj3AF0pBYoLcwqjsr93VMOSayoSZ9x8qte4loJkzS9bgOGzlGHO3epM9zQXd1Ge
TUwvqI3V1ttcE1OjMlKeDE+aFeduRmVwcNHLgEqOhvTcVZ4Ms/Od73/D3xTtGvWSdUlGQgUwhotM
7R8p0z9IFhPRdo3vDUXYeJ6SNlYZ7YsOkO3dGwEmUwwTfU00VFZZxfo8NDxET+TXrFi5AADw+tLj
7hqMwS/meTY7j0c7b4W9mkmDSp82Ict30ofEAjq9E99SB2h4ky2YzcTbRNxIGSRixqKbrqf8kEvh
rCUMePGVjnEeCzItwYygxyjCNIRG+gRHS+sjh79shhMp/qsWQ1wF0lQeitBCqhomG5YE5KJlflzh
E0Lt1lHz6MCG0LlDgEnJTiC1DXw+8t2iTXyN0ZcQ0Mnn41ELzHQaLJc89sQi1DfsLXklgxYFFin9
wi2/lut9iUPHZGMeyHKiwBZ5yUAUtId7QLYSffX/LiVXQBSPZiC347mlCLGc7ICVdfRJ1taHP6ow
EClMA8pFemgV2HchtzihljBAtcSvSTkd909tlcKwXNHaD4S4bwLdkPpJ9GYZUjgJCzcSl2eFcwY6
so0+2Bqvi++10+cMOHhwNOZNwY3MmpD5PKMFm9yojhAC8yQVgcXS+Wj5xXY+vvfPZkcXyUoKQVU4
d58DEXktELO/QePBkXOPamvXwfzdWJVQqywjaCOXhAKUtOJBqGBQ6Ne0Wjq4ag/00BT67hh9zwjF
Aqe+cRCT/onlf021nWWibS3B0OS80Ap+4YAf31gSzYX0TR+bJ1zNs2AczC/9kyd3cXVBe+BqleZO
CMYdiaNP2z+VqJ0Tz4fphoNMEpP2R0g3Dcuhrw5rGZSKORJJleOJzz/r9KPEFyyQn81eOBBltvFR
1VpBmyHuEUGO6M8uKcdfNW4xRHaKsYuEPGUrXTFPgtp703uc0cmASqMXNstuKMGDMPQtdvanDX0N
rK2/hjOBGrkwp+yYBwtzVvgM0aJ/Q3W2aj1EhsZG7/f/qPOaWqez4dx2rDLiPEItmZ78BI7u2sbf
dMUCOeW81Dg04hTGyeX982Qo6jw3zLNCJUpVKkxCFnopkgLQp4OmwAre70heFUSH4WE8s5BQmqBA
g3UyKKreoyxsuG8mQAfJe9R0JMfTjSlX7g5BzxftcVQmPqmrk9adIEFRlPvCKypnJrSgVEOD0Po8
lJRrg/UwPgrvZhKrumD+GCNU6aMWT+QQ6oOGnxDk/Q41sy43bal0+8tS5fr/wlStBnUjM37m1vCy
o2JFwriYL5z2J6aM35z2dN31OQZ0QNzsFp1Qp4CsJJZwY7CepUzwP/qbYYTzgUvmmUm13G/++W0w
IOc2nxlFvaILtmR6wfOCK2Yvlwn4rCQmAgTbnxbP0GavN2cbkLemuxc0RbsLlp3+V6lyy+9gFdg5
5BYTCaycJylcydW4/lF3kGUxhlr3TGYenypiAM/ME5otXMvrXbrVKQh5z+8RnoX+OjCvpUx6DgoQ
KwNcBTeon4c0TCiFe9/EkQZdnRkKHdtghZ0GpPqb91MJAZlxileT2C6/psc9wJIC/e8wap7aReM9
SCNZzoUNXWo5/h7mXF0qEX/4FWcIqCVPPXsfd4pGL6puvIxeRX3gy/Vo1A3KbFYpf8lKCN/4n+Vr
TF+gA8Ws7u1t+Gl8Xcp70LsDZ7v+w1EQKROTEpNkFOiLaeLeF8WbCcfKdtHlso3J9ORr0zmMs00Z
QY9IkTEXSLQSTmw0+lYblydbDx+tQRM4/XIYe3oTte09+wk+8FC9y5LJluyWPHDGOXMvgQZ4RybE
8GOvaG0kYDue6BwHKLQfOoonVEvyIMD0xrCY9ovf3yAZvBS9LhVOvTx9eCf4DmFrBYqw+Xgg7Gj+
QmjtaX76Ze/byCBx39i/VpqFfTcVcul8xoyzRO7Q9ce3exnSKz56QTVydhNbseq86pg/1KtDHyjb
jP7erUCgnabTrAohua2r7vUS2doz/ExdZNZ3C+nqhop5i5XR3q0cvNWz5Bj6T4JqSGVTStZV+mvR
7oLd4s2Xvxgruqu0iniS5NqWJRQrdy1TExT5uVsu3VFDsfY1BTPE+lSyZpHnCPUjTsnBIFojOwbE
85kyLki9m9SQJeyCIKo98qK4lzlss55qxdq3HwNvyDyjDMXz0oqUP6Pwjjk/UDIy/4dL+da9V/q4
zVsqTQ9enzUbZWc8reHmwhduiiqVU+bXaRcK6nsBwYM/l4pjcsSKluT4x6govN/RgoFKO5MF5x25
APbXdd0FkqMMrGD0vQ/FS7F7y9QQjP0oigAmDgNsKHayxt48xd0HrRtmqK58G8mFLi4cJ8NlrJ5d
fsuqoY6hO7SpImB4wPCNQlXm2TG699GS6rdbf0OBbCowT2hVJPJP9XFLfEIY5IZs/Bu3lbZf4/H9
cuAam03ktRpECwSJXuTDQxidj1TYrsSlq71vhfoD7vEJad7pb2Ez/PQNhvSLz3RgNKt5llFkRgRS
XLYAiHS6eraG0qWMJXMvUNG4CxXBCKr94vtsRz0lOs3f5YkyeKYBKGAdMYMht+30KVzyQDylkneO
YFuQF+I+VjFU1EmwL5BLbb7uYoFdT6o0hNe4AdDaCRay1bDXdfon0Ofr+HvIo+BGWKdTbuJxWRp6
LtlMbirKgv4pgthjkqXcDIx937QnCc3SLlg+rlt97psdeCu5vlopVlus3a4FtsBd+7Ro5YtP/jGB
nKeCY40U30rlhxpNqbm2C2DRCB3Ob/bdW0xn/S9BD6c/x++Ou4yp3RIgD+zVaY3GRIcuMDIEU3jt
duJNxMsoto9oJ6c7+RtwCF5J/hnXvoi8QAskBXYoc6hSimF9x/AT9cxtuapS9fl4NKMO4bbj3bwz
MuHIeXd/3T0IU0bZVgUjAemGPM1cckeC3Q2fd9B96KunKQoXsjmcr/TRoab/3XLEIzs85wVDnEzC
rM1GqxtV6B2GXy8wOylKzNUpziZnYX0Dqh1N4ePQg4DXt3A56R8dVl8jeouE5YyinmL1gUkGa2rk
pPeKvxgAegCiUpVpaj2yQ2mv+cVxVUo5d5G4RhfAT89XpFE7BrTsuXvxDh67xji+SkYjngJqPHP/
vavD9qXJJb6CRvr3PZVLzNKioMacyV2R/qCCm3F0n1PLchDngV3YTSD1QQDDGoIyvDlpJjASXtLa
uu0c+IDr91Fpo3yxRsskPj5CnoX7UgY9nomoWXdl2FVHvR1Wqpev1kKBwklTAAzleKJ1rUCSPMI2
HjCIyRgVrP1Cmz6vb7adR/56gFEMEmcMwN4Pzty4E2gijaRECBrkpX8/eIz5SU6pImMDvM4jEdoO
t1j7lfvq83/uGIx9gn9m6hGfGxKLHLoBieTjF05ImS48J3ac5K5rBTev+zIxn9iuY1gXUV5Bxe/L
24kCrv4eYXTNblt+kwl19kdu6K46Tdv+DjZqZgxRJWB19437BekUBY+AZHN5XnkOyTTmqxlJOhuG
CpxT4+BK5rARqwbopFgbM3J3w+XEC6OTBRSObzZd1vqEaNs8PLVlkNoSgKCPqAp45FTuT33WMB1b
bwbhBPds5WQ8wSWOL59yplKu3WPAmiZGfN1zHgOlQdqlGjskcYZpCU69j7uwYeK5PmO3LRapb8YL
f+gx4ggvFkq2ptFlpApAwbUhYeS8Nmxj5QQWeHgYC/sG5IGc9nq0M9z78hNU3nzPYnY9ZTq+0RAl
mhQgec3tJeL/ii9rD9Vm6L9ftnflWyayL+jpyirZEVwks1d2z9tuIe8G2PVIMA7ufMQjvX0QrEVf
RptQM3RTmGRhL23vhOx+cJstgOrUDQNSs/A9KuokBKHOeyThW1ZulImZsFJDFIvkoy+81h0iAxMu
dDsDIRpNQC/CvGQZjUN4+Eo3bXIQIWjUcOUxZXIr7MjaMNMN6FggpiCWItk6l2sRr1LZGNIp88ci
bbTU/lQtPG9tsxpB3Z3+XwxHRcRmYq7idWbds6jCeEqH9gbBu5eh2rco96khmKbrAY0/dM2Zvy+D
6euiJ4mTYLkkJ3/aW8ClTwU37gHmk1jRmmhIM7Cf8gAz2HMdg9+CuZqgQ4LTnNbU6aNFJMUsvIL2
q7KTT2hMCOsfEn92svDAhEpebZ1cJwuC/kUW9yYk0DhCGJYFY7MW1zCK7SwFsX+AWxbttwBZd5TX
2Rcg7e8WDAabYKg6pinyGUdJFYS+psH32EUwQJu4cFbOVRNdVBGk1JN6X14P9hsmThQb7SD4E8Py
lmgoZTMC9GXwrbcGo34MCO1n2QnMvddD5gUlo4BXvujpct+r/CgNz3QzGtQsKNG9XDgBzr1dXbK5
73MCEXua1HaTb3fyramquLEjEU0urpDetfGb5OB9a97wCdHRP1X+JQ7vqk/2Hs1cE7f30a3d8npK
12xa+xbGDHO45juBf9bMuVvt55IgAwAFxXAnZRRoOS/o8zeEJGfgINJSo/eJTEFgx7pfJuP4T7zp
uiSbWWFmdBF7t/+FpA2W1BJOAcce669insZkutNGHrT+7F8KieFKx7KYt01tC+FHqQNknFZ6hCo8
YIq3/vHjLjGTUKaaXuji6IZ+yEcNNoJb2IPBfaKGT4uUD3xCxOyJ5mniZlH+usBFfUJvkTkcCDxV
r2CzfnTMiXL3hiYShKLyqRthGxJagPDqiC54ByXeVbPa4vtpwCwUW9D8GzB32usZ4/MmXlTI1NHJ
W/Lrbn5R/4xPctnMFR+Q4efHTgOni41qL74asJsJyWDck34VMOLPDmj7bpR/PSXf5dU8Mk683j8A
yzN2b+/ZZjUCnso+/ntkXYoEQSMcLg69E2UYCPuzQZpcPknw6SgjvP8JscfiZdUNxRmT8ldCiTdn
E4gxM80oLEYXogT+rG5cb7SJitLlnNPSrbtAUbt4FCIicFsB8TJ9dhQf93wd8FRYYENxYq51BSmd
UuagMtsSl/KJ2XB7iKAY5EOD3d+EHXJcbwpPybhW2O+BOl3MntVz8A8e+bfXKLzMAJcdIjv9O8i+
Px8d0McX8u/u2YryRP1qDXz9/7PBjVkfBYGOQF+8koPnv8b9hhl5H2Pk5cPdR3+G4C/23TH+PnRi
q3RKg77D4TwoSGAAqNO9Sr35PifFD2Jr4aKtGzajFNIdvGQ/GXQExntEc/5DT7CKj1ZQmZCntQP7
GF5eNsKtn6gU+D2iOFTGrL937W3oQbq/Z6jDKKWWdT1FGQ1GUiSWUCKcD1eQ/ew1qmiUYwDPC/Tk
UjztxtuBCb08K+hgh+PdaTr4IOr935X8a3pusHtxm4uvqm1BgRwUOqnFiY5KtB2sXR+7hMpI8iVQ
l1m3K6A4oAxaUJa0UwQf+MD00UPIu/rolLEQ5TZCmfW4gwuQUVq6bf3Cyc2St4yfcC4qD/ZbjVb8
aR9LDsjE9r8OCPSpXOC5srXtDLLcXHr2IyJ8LHOoA10bZLzqh6InUsC9CnX5kvpT3xeRhR+UnYOy
DGVWJCKOA7SCcaR1XBN5hlDm55VSJRVED97ESvlWyBFglWFuzsC7RFFOQS91hyzQGf5ISX82z8eK
Xgx8Ed+XdO2NoHCnZ5N4mKKtkY4VechZ7Bv2+8YsgI8HfRJPOVw3GJYFqw7iGz107F3c7Fahi8p4
S9lKN6fqF0UWHoNnrWsNVlkjgDGxP9gqBXp7Lr6Q1jX1Bz8jazatVBrDikVTKAd/Cd7Kf5m6c/Nf
mDCOK6R2M6Qq5lelCL1M1i8TJbC8ckky+WZ0RVw9kDwHvR+D/eWnVBidaaar+xcJhu6ZD/uK1Smk
hmEyWVnJgrpIiwg7+4+cfnOZ3UBfC5fagmpCXSemMPhVxZgd2yoNOPSmWI0wr6bHNEJI23+BvH1+
Q+AF9zJAHnoYHrjGuvXZpm0LHLzObcKFLCK7IGwUckXXtM+TofxqBERprsPCCg5KUx9LAu9u2Vr/
eoYWVXgGEr/DV9OYqP/60F76rndxcdmRYpNNfzVoLU3/pzzHH/WC90yM4pR+U7z2BKjyl0qDQiiC
Ja4e3hKQH4eE/wryUEaR6Bg6OVnFzaGcSJ6r4ewGWXaaXkMyeNVHcmj3MOh/WHKQBPN2moKLLn7N
uk8gQk2qZXhHevJvAlxro4kCQ5p/9WtgoM7mmhTcKAxfe9fnAH85U2Y6m/JwN8B34fl4tBTduuoE
Kt6H+WbEzzaQypSom9tXtCnCNrr3DEPtspKD5sU8UmcPjo8TIxiIzBDv7y5rjFLGAJgc5iDMDsfB
X5mOYKq+pJpNZ7PengTeNWm58uZnKm+QruSJVj3VlUUd5Lrj7A9NymVHkPCc4dre8FOunvPVtG/j
60XNnQZ8a96+77KlLjwUUoBhw7GVR9e4FhFttQuftqDfBkmPmqeVi6FJiWx3SsGCj7Ai6nmdkm4+
I/JmZEnzaiNzZWxz78fGyA1cL+ihlOei8243fh4WHv0ucXcs/zkX750MugKLzu5WMRpA7TN+C9Ak
0AU2Q15dmncVZf7sWDjHeZj9jYBxTYKtX5TwHteAEZNhDgrH1oT2RJnQ/x0O+w0X4oCirtCyh0zU
kY+z+5SIP/WicDp6DrnWLC34mGb6MA5Pqhk09kzpiA+NqwuR5IjAGS8TL0Yt8XSBkMFDs9pbFdoq
oewxvnzpu38djkenVRQBfHu/Z8BNpBDhqSPzdO39mNNItFnlJ+F1P6GUm/ctUGln3udC1SgHS0jG
Rofa4OY1vivz02WUmO0h1kqTRxr7sQcpGsu8wJ75L09YM6cT3n9dj22SGKOyiRbvJkG+5w9Gb1cg
KAdMpcWFc7FQfkIx5c0yqaD/l58ibUWTNR/HDlzl7yosILgkGLmWIR+8o0958TLuY5j6qeQzGyBj
VjzIlbCHDRkobu1kt74FQc+6esECafJKi9xjkxs5XIPk/j4i5ageSZsv2/vtxSWlIkPj8PM22OvQ
Z2ZiNcvYlkDTNE8RbzgVtrc26kFV0AW29YLTzgOgR9bCFF3+rr37PgqBQqUN39YrA+ijLp1Lnotj
1q3c45Y6qCigAxY4xjJGTNofr+dmZHn1gXP5FTiVWa6SyOtRKkcgmapTHinx/+ah3arZqjRurG8C
w2K16VkaFMFHB4jCbjBVoN/9unKqWwNrF/zkQvLa7BGqRhZMC8wWgdGZl2qaK/Py+Q1OorSZG9BT
D88uXBFOUd/UL1knmAFXXB5blU9aFeWPa5fmo1ZUuaCAyzFUx5Chg7AM9h0BYqAydCK0MaAdk1PN
r3vKtiYX4Op3wh41RVxv50VadAiqDnY06DGnQoxJDkSF348Tflar4Y/VGutxR2KCTpAWcha8+sHZ
cTuizpbNE/sSoCdAJsl/hqdorc9+NLKEoaR/SNgpSDziaM97DXK2raLL6xe7NunhKKKafINnhBgp
Gifuw03pnnLpyO6LTQoh5sjDJP5djxwH+oIzT7zq7tDZuocEwAs8IN3V/sUhu099aU+JaAgHFshK
hwo5j/ltVV6btNxjMX2XUMBkP8ZDWQ8OvDsTN+qrgmF5gDdm2WjMw/zeJBjSOT4VZuYM8jtJ2xBp
7VDso2S34Jk678efVSIdKp2mgQJi+TfNZTUahwI2/RhhsE9eu3ix/liKY6Tzva8DGow00FkAsBlo
KSh4qfbOMX5fg3guTsx6zz36ADp9Y68U0/HeohYVziKJNfPe5wZ1qvgunfRPRR4lv85JxecyU0Tg
XDItXq420tb3TotTQaqAnY244eNSMU98GiAHJ1BZoDaV8R13sjwEq1bOepESmd5ti8ScazQ8DgiK
kLQjH9a2yvesnFnmkIch6ByKrGVu+CWa0c675F3jz7Y1cEKdl8sNhKoJ0itK3231awvprRjMd2Di
p4AjsWENYgRNNTDe5uAdQewqecNzq0B/VXzYRGN7mDeawf9Mav6ZK+5j0JuI9doL0Wi+UgY9AWvZ
Us531GF8NHEyi2NUC8WnreDqka2Cry3oBkmW1TvGYd+ImJFhREzWFldi43yyeQ4OnHCxwkO6KsRp
A5f+5PQQWsTrGPduAlvomzjiM4TpAzFr24yZhkRJ9P3aRbeLoxJIPnMp8G6/5O92D6KT4CuigaJT
nuv72710j8miSl3Hnj0W4i5O7yDKi3PqyQo5yOa8qI7AuDf+5jJPW95ydxCTmAknhWivDyvbrMWE
gsLVJnuRfQFXLQDKH52cKCstFfjD1IFPKIdMmpIOMxZGvUWfirxXEtud6j8JYdsg50uuAhqqxcDw
wL4yNvkAne2ulRo1sx8oTBIYlC28lMmXtrP+KMGWxbBXIabbMYXK6ka5pjSrEssNHReJe7jZ8ZiS
BN06tjf+2iXhNRabMvPOP+EVx9qu6hWLng4A5uEK//D/6VnD56sK2pUo18PjpdjvdUTwEFVUUsvs
qZJ++YYwpzFZ963xs6iQMqtRiTTIT37dW+yurhBZXMzDlhWsRR4n++2chced3xCKkqV/2EQ5lGeL
Dn5zTSk79nI7dziSN1MA+F6+HgzozeNyDOkrtysx4wZ3IPE1RcYbE+YE/PSXSVGNtCkeT0n3UF4F
ydqh+ODoRQEKiTomLrG/BUfdUcMhRyc1cOiRDyCH+Xrg92NkXttfT7KOERBpnrFU7SLErCBRPlqI
kBBHZkJkaqyTLTC6YrI7J0VCx9QvqExicYqKo3AODwN1OZWFvzfLXAuQWSNhuqHW0E0p2F0FTMc9
h266L3BShSnJWFU8Vbw7SxVKA6H4yutl7U/Qr1gWRRDx9dPFNhLwme2mQ7tNC/UXDo2N/RaemDaW
xfuxY80979rWD5yJotrEipXCJBN0MX7hxGxE8cYbrCE2G2C3FQBxDqtLwafbLNrCOqEl5yw2hJGI
x6E0dbsg1UrxUUZ5krfnP39f0YtYwqNWmQ8uWzWTWnmghd1yIC7FGWgMXpVwKXUlY3/TruLIJUmc
Q9KoFu/MYJK2xu95tj2DouP1B9k65EU84u2hgyeJjUqHJD7DZm7vImRfjdgv0OTO0CnY+P+4tJs/
uOM435uxJw071vpgUEQa97hYrcoOC9JXlGKnoaBPPSf6b/oJReXs89YpSxPOj4imFWp/rA/85DjS
dTQh9/Gf7iLnjFwpVCUIusR49Dwmee+d0z4lH4C0HAQ5ONIR3rBu3RtDSA3YteY+B/MG7kCVuZkp
CrJcQ7uNKZ5tU3d4tKsd9zlzUFEHDp9C5fmcTzIMZOz0xIbgySlF6ntcJ35AtuydnF62xFY+6JGs
GvPytfZCd2xenFMAoNHQkxKTIjLYByUdhL4CiF5lRwcFGhnfR9fi+HIc6PXqX66Rl2rgPXjY8x15
pgpQ7WVjrlg8iVndY5oNSQStA1OXmAaDVkI5eGJmK0KIO3qDjz+gSkWcmKe0QYIhl2Ya2SlDQW9J
m40m7iSsu5K8BsDRECt5Tn61GmlT1NI7qjXQXO/Cy4A9dWtICJpZqoMI2hEQavPKKqJJyXQ4scix
dJmd8enLwxNjh1lfCEZLPeNNmg59sGmqHOW9CzIuEqaKspww0tslGkkG21zxmSm8v6/TuKmIACB2
q1my6W4m2hTmB/ieKd+vTdLBGMkf5bkhiXJNafx5ZQyoq7O7MBOb2ZRka5bLcY0Qh3ramlmpiaLR
GXVvSHVeqEwCj1Ggl4H/lk3YKzmv7GHXTJaJ8lnz36rw73VqxozWqWmGo+tP0ZdUEY+WdNhRjXQc
4e6iAPGwDXw5Yl4NFFcB0IkL2aIV6/KNhQ9vovMBjg+1loW3hZbjmCB/YkbX+Vw9lav55iQsCptq
OAwnhpRCQ6qfDgvcsbkEpYSwMsDo5Z+FOf904OaTI6+8pRyxdifIym53suHLzq+XIq4gScvZSI9r
j/3TrZS7mTXv7vrsUbjq9hXe1OqGgG4gxFEBspsYa7V9E39oOjvy+9onC/kGjWxzoVZ+yrkit7RW
xv02HqVZyasJefnnYBpGN5sKtKGkMAlAetEVFQv6YaUJ5KIKNT1Uhx/3on9Hqav5Bpfo79PeHYHN
vmQPattHvw2K3TDFYkM10KJyUjk0F+XCm8oEvq6TsU65Irx745j0WkpmMl0K3iJ0uvvLO0mrCKFs
BWqjUmF3azsGNqni6YtgX6BKTiK1INXK2l3RRPL5iGZtaLZ6sqSS2K8o4eiMPmHA47VvwU1IulG4
LyCStvsVCYjTLFJeWZ9keqrrcwv3UPj2AAe71sydZw2zPdKKaO/E14fIJ180hljdZlFE+U2Dmekd
NTD6XHLp1UgTMHj3R5ICbNgie7PH/T9EJJsztD/yxyLoasrXbIm6vAXVouXLtbWVfltI0c++yF7w
4urwM+d3eEyLwGX6qqZm1qb/RRT6gxp+Yt4EeGIX67O4fLSIL9yjSFDLOwTikLOac579egmuDhOJ
8/khrvNeBaIGahYUwUoNOBP9Il6DW5B7sqhFPibeUlD7VPBYTcmGUovH6pJj5pBI0pcMYr6/PMNl
mUJ3VnlosRTBhZ6/BOamvtO94ClcRJHp3wl8k+w9ord3CvDV9wLiy5tBBytZL8HoDyADBzKNxIoy
jqNtUoXYXFCkoFLrOC8MIeA8RddFAGWZ+Xl9zeHKIKtuGQbY/tMtVchHapULXz3z96bBmKdgRI82
+QSGL+qXyGOivKQ48pF/bLDZuTvuaZ8kuXfdnK46zCvS0+9iyUgLzL3jBq4zwd2BCErhG9/pr5i5
PLnRwtoDVgp1u1ZtjzLaeuHQ4mIpcIeacXuol+D4l+G+lIvg6i6ptEUlupq2LflQAgberx1fmUe/
rFG4CgbHtPdIDU1P+rtB6aAKAMsJCwyiLELQ9QBypgAgXtBZ66iNidc0amv0RNVCZJRyhLevnM41
g9IhXFMvkc0ESh92+4RkRAW4zs5M3ZwhAoYeDbQ7XAfu7PXwLHhK7j4xLV7GfJ2CaK9hlp02nppM
5zEfjzy8U705gDIHJ5npqTytbZVNud46cNm2CMN6keNR+UEPgQeSjh7PxxQnCDR4/b0ghFLXVq9O
KYe6QLxjIZMMZAhLPnAmWvRJpt8KhL2SxJKWgVx4yctd3+/i/yxGg2qiF/XP6vx4jjyO8IHa+Fx5
fg+BgI41DdcAXPG60nrxKl6IfXYuggK0OfQ5WNbcMpOq/rVvnLP6AiAupVA5yx4cVS46viJtEhc9
wDHQSd9JlG/h7rrR/CQpVp4KvJFHuuLnTyRJgpCHB1Qrcia8XA6RVlcEl64Q77I0EE6JEdkGBsjM
MsUc5AsYMGCtH6K19k20aY8tTvrlNBrZCDMEuOCXHyK9hhz8CWmns7nTPHi/6LsJS9TEvfc0Xm1V
U9B208NBdwTs036hH6+pukI0RdvP6EWZxJEA1pZywh84R/vgUBI5uar0ao0YElovRMJ/OaLO6QM9
XD2xfyKxzLRvQ8O99D8HeXYSCm3LQfTNwt+SZX+Z48dsiNeRuhTti9h7/g/oX+xBv3TyGdpw0ofy
2VX6ntf9W3SGJzUcmmY/fcXajRcLMOYJGclI99/yFArFLoBQfzxVqIZLIM3wo3x7OEMwoD9rk8ol
63V9If0BpUmsm4JzOTZIidhW4Mc4eel3DIZrWINLa9yuRynpz4ks7RsdDlKra8XoVlmHGL9E/jkG
mwWEsyM1UGLHJMVnRZ5BnqQmSrZL+naIVc9ICMXV9/rb0SLnYr/CJcKkAjbiye9woEvEiP8Z7Qa5
teLTVOXheC4hFJnt9HnUI2gaJLB7iH7qUBL/WKLm0T4laA1NHp6j1UtJxM4TQL9LizDcEwftBfUJ
nPQ7ERwFZf7AbUmUCNI9QU78ujmiuyUV0yTIn92qjEAkGMm7Peby7AbPvNZs14qvkxHpOh2yM70T
ttagKHIMYXrYSxg8rbbXQb0yIdVZZcILZbFbOJzLUzCW20ImataStr/IUcezqcJHX98hhgHgzIWP
GjXrKh9RnMj8O0y5dpFgCt8jkX/wf31TGZMyXtx5AX/iuijCteTGIGyatRFdvn0zvA3x4W0bxseX
H+KlidYSGb7aKg6JQsxK2OiSmeu+lfgFHAN3k879ioSKyI/LvjsR5OXoidQ1wtjRUmDMp72YXWFE
w5v5tUnvxqBh2B2iJMSQYiH/3E+Y5VIKQr9GX2AQkKIEuM0BSQDJ/M0OQMWIlIN5P32G8wTrkxvr
qVlKRzPnJaQxCldNNEhnutBEfhUou0LEktffTjE3IZvgS7Z2CfftDifFZfk1iAxCtfAzqboDlyb8
RAgrKaED1heyjN3nt82QzuJyJVMyWFWxnEqsrYt0tGxO5UCzP38/81sftgvBH8rh1pnUXx4SF5Tv
OGwsvsj53KnznaLJV93yNG46eAbtC14pB6LcU0ED+tuC0i8XrfjceX43mtxjhWXEiJ3xCEEnZVZe
EPU0GOwFQTbOt0kVCgDlXyM4fC11LwaBp6dcfYMENK3erg7KD7GW9wuB9/+uYr/gn17FF/zASnA4
7OlYCf9GmuauTM9+EzxiYjSPcROwafRZLiPcTQ7173u9lWjlXXmVkXeYqzHc/3bEIn1n4A29IC16
m6gw0CyRGZ7mKQO0UsxMHtPh7m3lBRNr4FUBfS81iPciKNnPQ3vmI9xBj2kyVXLNqWkF15eQNfRC
g7o5e9g6tv8jNJQHt+f27rGXTR2RXOvfTImrySGchB36LVlQ2yyr7iY9BcPMFDKiWzxIuhOZ1mOg
FvolMp7ZoF1re50GEdJ2ECM4iMQwDEzu1gYcDnK5foXfhpz5KCmp53mrPyWlUJnRAO2R/Ni8+vvU
YfHWALI0i1EAl9u/L7QYp5mtNC2sMCJcTyYNK5t6gEogm4YcLvdVN5hQwjtOPBX+W+9DOLGKy8KB
Go/A7+y6icD53avH6enHi0aFIuOcm5gi0cxS7hysPgGBtRBzIuuzVWZB64HVcHLkjeByamNbrB6p
+y2EQr65jYDqtYpr8JevSNg3GbP5zHb+CkBaAkHsFFZ2UHoqUZd6dpLdqR5hw1/YwqCvX6lqdmGc
AGQwAVCXOIP+b/ZGTKiJZg2kM5HYz6qMYDagVFpu221ggk0CtNgEGRkv6H/yoT1TbBzsm++pzOCw
Mxiid1fY05ZrGX706SC4vomF408Nupvw6qiUhB3s381e+IRk+iSrUDH9fd8vjJeWv0XdTl8Sn0dB
cKqrg5rudmWvTIYyeCKvwhIXc1vkua2ukg/14UREZbIXJ+beKiAa6rlc66/KFgUM0qOjTTdvcxhg
spbujgtn0DKGUptDBM+I0wGDVAaigUorCLkIkQkmeHgimLZ6ZKVdnA7ki5+Tc0WdsYcf2MSWmdVy
7ZDwMP7tuv6/IgSX/UGlNzKVdLJ4r7hVyKBu2jY9luntq1m8lMZTILR9RIfnRr6GIsY6311IeTUu
1es6ZJtNJzx5gCDuqHI0hImCprfv8SQsKg5kw1a55PftIqASpX8ZH5nbrpiiOTn8yi9fWQ9bN+r2
qRRRGGiRMV2vyGZ8Ej9o9qWz4RPR5vChNVIXqe1zgQq0XK3Xs2MT7PYMqSJGK3p7wwf0U9ob06DW
QCm0f3Z6uTqUH4CS7BYL88gxsJLV7Z55MwK6FV8/ipd/89vQBRpYwlkvRiZmCc91cPabDBL0Dvm+
Tcl1OgJ1JuKnNfoobq4vfw68+X71vmlEP84wVJPrBaseZW0/2E2GM2w6ed9bg5aTVkYE3EYFKspe
iqulCB9TP+fDGhanN/CYNoLWFbA02ye3qmaO41kl9vlQIGpUizRKQlaeuIv3XPFeTuHYqQZloBZf
58RmjYTDN9DtJzhtA+svuAHyVOSIFh8OBtkUEdpJu4LBTmgeMz3UXrtk8Zxs1HiqnbPqCvEt87MK
OWPnppp4hPfAX8jv77+iaTDG3odz2s8PLmkLvvsbBBwK+n01PfyEgxpWc9CQdR/qMB2+YrOi+sKK
qwSnWbcg2MkuiIns6CiSJ8QBSP2gv796Ijz+SHhMYEPFcxmbeoGFh9GveEESYfu3ZagqYUhShpYC
Q762q+QggMomeGyJ6uD8/Mgi3QTaU0IvjVx93AlJ1vEuflyvipZu5dJ2SgR2KUaf+Y/5+pzNIVam
WxFDt9QaT2vTkQkwvm7SYJsYWjuYZ2PT8Rqp7MMGmJVtEV51bbSLQMyjHS9XUTaaLh4uWRnyX07g
wsYoVsyyc7H1Zisq5hN/aRjrLgyqZcuBIa36YLEH2m2YMk6K2BtNtxLN5598q1WHraGGCAKMmYSV
8qKUe/0Ls2mMS2Pt/WVqx/ufVKshQ7iCuOMrz7vq3YHh77n2SLLhNi2QRYgDTW4JrpEhr8qUFils
yp8i7kmvHeLkkIKJX89/dx2b/8npi3FrRzQOWp8M6uJZXwurTlrSK/nUjsr3UmMtbB1c3TA7BcFA
CQcZ+BFLvlcBlQCteu/en3gF1Wh4jM5TZfs8uySUGsLxy6FuQPDkpvIqn7eSUWsv3mnYOhgK2mkB
NiZPn8MmCDCZDZN3Vw3cA2nI35nUt6RN3GWRDiVbM7n1RVSUIU08EcS13zZ47R+gfZdvVHNoy6Gz
Wor+9JKU48DjTL3+q8hKWxLzx8LbM7qhFtEdGoBMKVogX28Fa6NZcsjvRI0nz23bP34mOePMg9I4
e2N+P9rBq9KT422uQ2jgXbWqKOZqinKExp+55/U+ZkblvIGBSVNhOeatmXat1ZnaH4LZzrGo7qkc
vvuh8UqOZuqiuI6lkQOT/yJa89cno2F20neEeccaF4LV1nwEmuNDrbY/1V4GGstDwkr2cmCi0vDa
0SkZ1/K61JCFH7K15UWJ1/jMUL3eOn4FftO+BsDECF+h7B7bHQo8hs+tIRL6WLwVYQVMRhlsrtZ6
XNME+r4KzxOcD7INge/YvwWTJtEOt7FoDgBkVntLm6s/HpXbgVu+cCspIhhKBqVPlXXSTRiG9R+c
WadPgxNAcINPFTo1kLiQgGryzgpBo0uWd18mQorJpeckKi8BtVAaKHnKXeWRPcDHncQMBb7nw4OB
My21Mhv8tqhG9cnviyL8qeLADszPdu5x3pHpWWDnYc88P0ipzhQ+VI1ybKOuNZOZuvhvcoQdcb8I
4E4UkEnPmgbITk6doo2Eor9l7X2Qajt3vDX93p8w/BsRluGuveDscKZPpdiUUZj+VTXyT/KmazFF
g74HPAOdUJUm9qdjYsHgXAGRDDa2nMjViPNd0AqdSFFVfBN1KjaWH2xqhxLO3v6h1fHBxc2fVWuT
2oRdoK+9JrfsH3yXQAZNM5IBP+wgeOFMB3g/2ZDbszynvGtMrxSzfEp8wYs14X5JuLiqzshHDgV2
v8sYyNjtu/+WIYIvyFYxLDP64oj8SICkbDfoyP8eccV63ujkr7Ma5TbYriaUArXoW35nSHFPwIsa
E8DwZlX9ynT+Y+53L7dFeLGQ1STancexuodZGr9SFTsiNVHOksGR71f7RqPQSI+oNi6A1IlHWc2z
ZKZovYN1/+fU01baZbF9JFFD7npG5SUeVxLOISJHqTGiCIKbo8JoQCeDdAmPYffXEQOAtHXgO7Iv
RkKEBZZMOHS3hi8w5aJ51+NgwGyPPCHTL9xPzF2d+SJw9YbbfJBAhoaQBl2nLH9F/sVui6kgg8H+
heb0N/nyoBoc7QZMfSmkUWZUfcZqYdVBkqNyPaMsY7CnHAzUZTMifXy+7WUwVit7FdoI/vb85kV3
CgKixaPYUQ237AOUZxfMk4vlZfUYXOhYesEKXapBGmR5Hh2WjwyBYJRU8ckxYscIyAKwVR6S1BMf
1CtKAGlFEl+42IhH5Ua04ct8khb6KyR94XypA53Ly0AK42fSVhTNWaEWkqRUErA2lwhKd001YFlk
S+fUHsV8Hxn2hN/BGjvSW+mNG/PQQ73GC9/0ZXiYZoUjNh6cp11XSEkfEtQOw+uDz4S7LorB4tMJ
nxREZtsi6QARnnFElS+xtKLAJKjljttZWsEcEidPX4HHO9KrM7l7eysFZhR2D3wpaGmD47ELHlrV
Xhnk4Ds42u3RpR93uzDKixVC5Dj6r/NBYpUgQvOomARzghtnHzp4lA78cij+5FATo2WuLQXtof9U
e8a0TTllaqFTdYaxOWPxQRVjuJuKp+q54oHfsOirn/E2Ki9A7p3jNRc1ONCdpK2uRVlWCBVVykA9
7xtZoHZzyA+aav1DROFvBxGYdSpe1CGYzu9XfFhuhXN5L3bQfTZUdDqCos9Q9iJh9yQGoVvRLcQg
lXidfmLn4UGZbdIZpyfXtk98Iu1dYGD6DbZ2EYrDFZc6yRnWxLlOBTZGxrdGjfazznynqFeMye+n
uQDNkfIW2N0HhWU5MaHENWEOunosUSbs+IM75QvNDqWnXQNua8Qaez4KaFR+acch4n0DqJSODtMH
U+22Apz6DnxUpD2szPzH2UxL/fmXGQKAaaVdKAZ4i8nVDhIR2WZDz3ilIi0YarwpfB0Ll310mZVk
RYOFfLgwj9wEoKWORfg4KrXeWtXFN0721wO3w7mlgk5S4YE924Oim1c6dDY+an3mKKGpSRIOs/Rk
YpaPHe6dAfvPhD2HFgfpi/C+/IJkAb6/31y1d46vtDE0N26jSoF5cmIMNSHLiW1bUKnjBa8ehU0z
qCVGCEY2cAX8wLz8171GyNu9BClY+vjEqqEMRRrxUWSNd34EHOyTYTFgnFhtkI/j8nVOrG+GDw24
pk21UFtyPpwjNI0ry+6JeCYyL7eNb1mrdM+1629B0pZ6U2pg+kn3C5Poy5orALOwV3heKncj86k9
2bPoBXTdvASd/zp2qAZGGIbrYa6o9a9QmW05E3dZ2T3PImmn9Epju7zf83/oUTVPh+A9ZQyhA25x
5hsgg11UPTOPwVJtWL6GCWQAh1J3Up+pfahFMBZSPbfsLVp9nsX/qXyTjMK47BmgbEMOGtjVxczw
dqXz8A4bDVT1blGkxCBagGbkqFx7zGlqbWk0ZVlj+iV54vOSfO6p5YNU9dE3nJBy5JgIuCKQBqem
iFJ7+QJQnL7PlKfFs5YDwo0DNV5awzLnedOo6arHxXiUm7Ep74r5JO2caganwZArSVp9kYl0jHyM
rPou34dPGr3fsIvu0wAeHeyaS1GZhrx+B03bCmsz9c8Qq1vApjqCGa8oc0ie4qrcHTQ0nie/9yV/
h6cE3443Eh47Gi6m+z6/kvEwhIzDSp8z578qyCltv5w/FcakwyWaYEmDIvjho3T9Tue9DVkrnkuf
RrippRJIdpdfpEgkMVVY0HLKMPDypK35ulmzUqzh79YAdrIc20GzIdIio3HgxEWQEKvePxNiUcyY
K7W26hEy5bUOVSn2rmEt7Aqwxi7+aooZ4ix8FnkkmoI952pCVyTU1k1U7NNXct6dBDhuDV84rXxC
HEMq92hU2Pm0IbK5ODNwzzNLCOWINDYfdIDg+2W4IUiV8mm5ack38y4u++rPL37bWflh7D0AxSfF
n3H8LKKUsxkBh/Q8Thh0U6U935PppZaJtPeT9kFwCdwK/RgrH+VjMwiDSlyV6o138/2Ra+cX78bT
k/DtMnwqf7wQmzyNwh3p6JeMXaCvlGJzfj+dZ0kXSLzhsKKNWWccn2BFD09khx3o5L96vnQU37Cp
vYgFOcTcI2H/lFBuGhpu2883czNAYoyH0PpD/1AN1QnuoRebJ7lEIMSyicFvjRXyOOR3PPbK//Fq
Tp2ilx290WR0LvgwH0qSKpe0XZ7v4Fo87wCQn6pj8hZ0ITBz/NlfiDiYNI88mMlp9cOGDbq4vLsu
sQpL3FtPNNuvR43bWCOF18tt/bhhZdBw3BQ2gDZ2gX4sjAym49CFbDn2nvZEaM/xL3biH4L5vAQM
L52Df8L6SyE0kpsqJKk0zUF6HujibbxMrbflYxG4d8W3caJhSDBIJ6uaxVg21ovjjaXLYyzKHhiu
GGGGEIHKA7vHXVehMmFi8txlZIBZtIRyKbZqbAx7Glw13jfdWi+pTOXPRfhtqp80BZddj5TsFd5A
rXhwcZTHfgp8oMygf9rcDjJvFnEjSsOqIf76Qp7HIsM5PYxnCmarr19nvxI4LJheHtptitCkOK5G
cHr/m2XYt9vBxvBxXz9wJ+4ArcEDmltXOY5mHIqEnZ1l3AxHvZX7zZ3XyaqP2A4wR/jBFDDQw5bO
9eNlETEcUegGIgQpP3YI1QD+2eNkd16TyeBOUXpKl9iODXbPkdP6Rxj3EkOGwGaJJBOOKQHs8LqN
PtDPnHYawllZCXEUeilA++hVq91Bwggcmra/DYuC1z7hqee/lwm6d7cjCJtT67nk/HPJcdh5Xw5C
yyAYav3DyUcoEotJwptUL1Ys0j4pQK4yeD4yg0dEjIm+vlkZnB+np1sFt8O9Xhu5QToFWbcsy1Nz
hUFr7Uar5+uQQaXN5HXnv+UYtTlYpqAY5YKNjATU0zId+C+mm5fu0WZCIZHWsTrCyxK7XXVOpDuF
uL0kQY63KhyVwwVdowLv7CMF6+XwYjfrg1Mt2aLQNiuP9+tERFGLFXkEdQpk3OWpN4nR3o8S6Eiu
6LEn2lL4TQHToJEoHLAAdEdHQK0Z6px04lBgRKy29m1STdB+P6pXjodfzsKSOVRdHuCP/W9KzC3/
ISTMjYUVFiXUbhFipFxxUBWn37/iZUEjaeVv/BabxnMRwDvUzaX7MCuXYJMitody/qd6yWy/V9//
MzlKm0eLmNMYMu0BiZ0hfkDe9PXUQjA1fwandMYxlFuwEPA644RhE0AkEZa5TK8vbWhzOTD6resZ
9J7SL/1Iay2v/J5zNIsMLfKXNeob+bskXixeWEKlnxUYYk2+eeJHKSfWSI+dEM26rNjagSr57jYY
ydW55Jnhh52cur4N0q0BJNvyUF/9NnYXG56pRdiTa68wN338/WHe29HdgFccHIezNzbTIGByNnSg
MuGXiAk00YHVUAnKNdz7e9/+qcN/ZQ3DeRGUje0syY8ne4HBqSk2r7b0gaPa6dP5cOAtCB0yXJU9
7+ZOLu2ZGxY4TnbPlGjHvL7oRObaT4QYWXWG9JMPJofzc6kyYJxAjtV1/IH5OWBZvZM8QEMjdi8K
Syy6DUlg6G9/yGpv21nBPyamdACEwi0AaUQH6fbM+ad8TfsZEwz+cd371r3CEjpUi3dJI66tnhIg
AjWXFgFRRjX4o0i6YSnDV6oRK8CqqTNnwzcK3fEdr5c8zCN+UElkUmkYBNl67w6yH09nyo/9VoCy
oM3iHt7zDUjRmo2pUEd5m0ZupCffLd0cZx9rv5YwCf7yhxxORiPNMuchGBduGdlx2noldMCOpsh9
DoohSLepdilvd7obxEC/pTR0/YCOrBvfJeASxfBL3aTA+CquLe+EelAPFy6lYkKBPpqZXraBMtN2
LeJf4EFzqc7yrV5SkGtSF2WdqjoEpquEaDImwoJfLFMLp06I3bJAgqbH2EaiinIRs3WdTTV2JP4p
IVOt+ps8+QcN/h1jjL77Nq0R6LuHUUiulAMGOIaiP2rq+GmQO379e+G4AXtWQ7Qe2McWFTfKVoKc
ivfuhtYtz/UP+28Pd7W3+73vxgbbuYidA0NIFfhbZ+qJa+vuBsVC5lzoEvqdzcw013KSqjtnNCsw
vm0dpJQjRjIPNnWCU4KfwDHFfWCLYw7EE37cAeR1uGzv1L7vf4iYmz1ICZq1VJCIVIFP4ggH/UyB
Ee4J+qpnjmaLlviWoAVOBzqRzS73duB9zQ5vOTUTftnhPlCvjg8lG+VqETjRqntxu12FQBfsGZdQ
EgnpWrXJ1rC+7zeFhlgB4nGhxNJCruBvpr1gKOReXnLVdOdMwIMdeYCrit3x2be6lavjoWkMRvf+
D+Fwk283p/y54fo4QvdidaX8xya9oPdG9m+PXRIDeHT9OPjUaONCZ8d4XKHumlH5LLZVkstOtTk5
YfUEg4trqbFDsAP1QW5ejb+GXZ5h6X7tSekATwqDOpz5FXtIfy+kWjnWnTLDoyeH0AACrzSc5dZy
RRIFUNq0A5wQBc3veas3V/Ka9qHmXaXBs6zhPsu/NxqecRFn4yv5hPPBSakywDvAITUWIMNsGu1b
7i2HKNkMllTmJl4lOv5DnHLFQmA4xRZucP7ANRzpwi+OshDzsDKouuGyv+BgZ4zJPzQBDC6BayA2
J81jVhqAxcsX6fGQMdMNODpxHrVPMLNFrxDHK+X7uhjzikIL7hpynXiuoePZ2ZStsePBnc1VhFij
ykZbEQJ+paxna2chP2SGujv0nxsJ9n5+WuExvxrdKUyOzaF80PCINvGE35rAjMi+hZJrXr35U+DN
xxcJxqKvbPWodfH68qpG8J0gaWVc1l8qsmj/FYCErp/+0EItaHyTQqubKc88TGKfHtEcbzFPwNpg
KJHAKRoNBEZF9wRzXCZ6MLCsTd7OrNq0hf6MFvWrIlXlfelyIoduhEWiqKXc4fuVsUwgKB3nLhQf
qobvtUN+17sRuxL5wuzzOF2sn+X4sG9vM9RGoh1RGKJPjdk75iwl1yr1l2IdW8lKRM0LVa674gcE
1QZGrCDyltE76iRZ4vaVq1v8X3l19/GkZ4l03nc+FJfyR6zfY9OlHgG8VLC3nSPZoiZ+u6806G/M
01EbWkSXMYzXfCB2oL4fAges1tvOSacrd3RcQ5iA0+FMhITemxWuuSjinL3ohg5kCG+Ouk3wWn4a
K+rFwcbJOGfRQVyoDLxP2fOpLE3TyhwQ9zkYW+gA1KOdeMel0vWNo/DT7IbBw0UNEOUhw3UaRZBb
RnyEYAJAcAQ84g1xH8TuABX9T3rBRrdOo9cqAzBRuvVQCRb4mMr99p7RCzLv/GcAdCMTCZc8scQM
1OcFaNiF2tmUxy1ggi6hmlTopbknaWxf69Pkfxnk4IeCu5txd/LU6pTJm8VqEcitWSSzFasFUmdq
PQHiWqDINd4/FKHg2e+fbEwG4evc0EgaoTEWNCvOECv9uPrGlOXMpfYScKNzEbkwVympW5jaU271
wMTDSGlHMBjVWDkUGBWr+dYS8sRSh8MWt91+ox92cLWzq5ffyKjtF5UnD4/g4SHTAiFK5T0XXxu/
MM4aDqN9h/AcxK1UmCF6ClfBAxAKaMjtYADqMFstwLEfNrDls0rNm8qMtbbkf3eAyuxgpTKte0UD
LawRJx/+2SWLcL9Lbq9e7fw2DApI8nIhcKImYUy1saDyGzZ8rNuZUrtLYMau108F2vfcVJkMlCO4
UL5smPLvKtl+S30KMRiyUgLz+E+7dBuQ6ap9/mpd/RcB54ZXQU4f+w8j7vSPg3vUCJj+dTsijDEH
B2vM/CUfEbXKhTZKpYg4RuMAsnLnxun8KCTcti08qLBZKVjATTt6OpAqgncYe8P1GPWQCGzp3sS5
41DBi+BhZGXUAXth6HojbxyyoGHUKwLXP/Zevc4udNkSf576HUwiPf1ZY7NOfv2WE++YF5+4JFmw
S7J1oXBDoiKp/DM67FLmGu49+PCxZqUeiNqBHczxH/Y39y5E8ZU9BW180ISxpoUOn5kJDzyIpcGy
F4sji4q25FAcSzXfKWIn3wy5GR8GU00lkAvVz/JMnajLjGSsYnJ7MLan1kcrDUIjiAiCD5olgTKp
EQVGmCE0X5xYSnb/CvePdGOtl8qKnyLF5UwNelpvo6gOarWXUyvGwZ25AhrOHBpgHSOi/PsNOs9T
72D/NZBAzJag/pzR5q26uetThe2DCUKV5bshnhZwXHWvWOwXI4HZXpd4Pr2S/lCpb2MEzcCItAwS
4BhDOZs2FWNLvfyxyYegdTcDbLZ90bknb6fG80/Q1a6ndp1lwNWMiNCKAPMrFeStCz/aL0eS++7l
laWaOiqv11BGT4aVp7pPP9jyuertmxJmOHD4Oe83/8Y0eG65U6H2RlExmhfCa8mfWZ4QelCPlzQh
EQtUELWlXLlp+csxXAOqYuzXc1jJiy/ASlIvtanKi+dpUnHFjdaykIQXDN7KfU+84U22tExdWQja
vIRXFQ1pmUwIQVnEy8+B4CQw4O6y0hc6zjuntf3GfaUX2n1MyjcrJ9IphbFyIDJ1dA0jERtEAiz6
uKB1LqXbDMBFMaFXrySjFOtk6dOx5wBiF6/X3KPlB6rlzCnEPEyDzBXHpGjP76uU49YtOunu/TYn
Rc6vjA+nU/8zaNaGT0tPuoQarSVFshnY15xaXY9gQBoGKYNrwP6vxMi5e+KoZ8aWW7DQ7TzNCAfb
/UEqKYPC/oOBSFbKaculJvCjv+BPEgKRXUfT7IRehORZq5TwnizBrPLgbCYa36y698zw4NtkwA7C
d2jFC8tphGw4fIuU74BIYfxljF8Uydh4N/bhcQIRfPgWMiE13nhzOj6Pwm+TsIlFIO4n6O58ArkA
m03+UxuJhE3lNtThiA81csPEtnrp9AfjvXmSq7f/EuWuCPHkUX60OxE0Wo798NnQY7w/SL86POFN
4LJ+WvB27xZSSbm5Q7iSVHK3LExCfgFbE8bU9OxbmxnsJr8gq8cO+o6veIv22JztyE+N5stYqQwP
KB4c+y1ibo9b9IkSSdNol/l9d6m2XgdOHNdl7wqZtTUY3AFy2z9wT049R4+481LOK0ervEvNkT6n
XsQ7jbpqfq6pi8A+gVJ2bO9Usjw9BnMo7Wd2LKbXQoWjGanYYUUscj3mcy9T4+RXPYacOhYIPSTJ
X+QMS7X0CDy3n8oeuT5Ct5BZOBoD/uA2KoZyPyN4akbb8BOmgLcCj433pTM2CD+mSboiGqRm5Pr3
puOdbb8dg2JMbNuvaLqB3Qf0pUKfUhqDKQNnCjMAvmyrhZcAlLzPMxyP/kHz1E8+z98l8twEfJS5
rp56jja3b39EMtLDRNfYFQM32Up+K7XDnZ/TsQj42uPK1VUNnwA78+AJmu20PUyjM9VWZ1vu5/Yg
S+J88MHAok3+Wty4KvUiGZedzKxc6O+djQAIE5WkBUo+pvcixYk3XpkkpciBjEHeRREsbKlZ/bKz
Wrfj0WD5RiKJyLD7YNA0KsKX6RVpSlqX1cycmOSEUj6zTDDZoDj1EJzFtPxROuX8YWx34QbQQrwf
Ad3d47axrJGKbs2/vnyfXt5X0aqgc3K9TW670uK2Ug+N6UK5OLzU27gaYY+qbpY29StpULi5MPmC
xUx1+u1No7cMkzZYtX+qDBx/z8vxNwnYpSXAlrV3ugDOEDx5MEIBS+LBH9xgN5nSqUmmSb6GsxHx
5W0Ma9XV+3ujP4wr/UkAPzrkj1eK+qu0CtjRTj02UmD6olbx5wslXVmEFySQTEmlCxG8xbsl4u1Q
fpk5sAoRi7sY1Jq7QQndutbBi6Owp3TktHytHe+vLvrcMQLPy6SpBYhQhaIDCJ5O7oufXfpZnNIX
Oi4JVsQGdZTX1ysPuDZ9ybNaJTxMeGNHhTx0rYigE5koHRc1VxBT6ds5sWGEeNLMSwfEMPycki8B
d7wwi3IpE5tNvcFMmsUYGRO3FAqrn+l77JpXcb7eRE4uDtKh+pY/PIhXwdW/GP5p/2A+b/owfrDG
ncMDcx3vGyrPwf1v69uuGq7BrjH99hsKL8/nBS18zbI7YNY2sZcnDbHMGx2pOaRL/siJkAfQDBm2
QpXMWK/G7F5+DGIvsdjrPg3ytXP/m1tNe63sB0CA1uGSiHNkWpXspeGFNzcvQv/8KIrp6J0qc3g5
MkNIGMJYzvYh0bJJyK4bhfOS5FcSAc5MpPx/WXcc/b8IfKoFJN+Ro95sziQddafuVcS50+y7Qj1B
m3c3Eqt3Qdv+xvLaSw3U+3LxctnphxaDo8Q1aJvwoLD4lqzxe2385KmKgD13EhNGzJLshDlmPiIq
x7d0UKx04oeflQyxfXj+bF2iuGP0VAnQGfr40x1uxZJVREtCfW9WRzVvOS+y7JYp59gByvtdkCVa
JJxR7mO5y+OpQsUdSjo8K9pSPMyk3aWP79A/YmPEaX+R0vdWIN++sZhCPAnuu+GDXFK7gMHCb4T9
N/m1IkhZPJpXlLgyx2vqrhPNLecYePssBpRcO0bzpzEUEGlPNreqhrMFI3ep8Bf1KhRRSUXit6p2
jRen4/CkSmgbK1UEZV2PQec5SHrEkU44cMR29AoSkSAUvJtg2NgDJA54yOx+rJrYv66CPIAhGqdn
QU1QoQJwF/2r3n41Y0Ljg95IRnE6eQsEnUFnPwbwJ2CJCQt3b9lUkAZanlQd1A8TXpqKgmP1EfQ9
sBZAX/uGA35VadWM7w0+RKW0dmkUJ3LQXbtMAt5lexFx17fRvIUkY19df6Vyj/DWk0i7t4jGBLlI
EPiyVb5D0wWY/nwnrg8AaXtYH83KAQnlI1jwOV8IORRaCa8QORr3/tQHZ1EARVcavo5IiKh/fTyP
usiJvYWvGIgYc1aKct11u2WjD0l/ubIZxKbTcRX9kyuoGkPUafhg1QMFq5IHZZqWRkfmbBhUHnc6
chNuzuiaNFpj7SLLhQ7vZTM2cN1VoeAG9YjHiCRAAS5kGmAPP5TRK6hJjachh1/l63r7h6c99d0g
4g5zlqBMXAMneC+GGIJFSUvF56OsAeXN/lQWvFmDpRvr0fLMyElS2byfiweapWev900uEsg6FLX8
7tcI2uWeALlnwJaF/R2lQYAzhvHRAx3qn7LzCMpe4mt8qhKfbWUNjcQS/jg0geH8GmvNdc7YnyRv
eOBM7EQOfpa8kUadtFnUVcV8Gcy7PENrVkY55srsJW9DosrGYNNkUG6fzfrDgJyeZ7MUg3kexWUA
Ejt72ZvrtYKCj2q3fkQfWBqHKK+TNaiH3UhSBAauL876nGnFOehLTO1A/6oMSWFsvzcNO3AdkvWW
5aXF74xeNvTJgIHGNCQAs9Vj9nbFQ9tixCgPpjfNaWdGOIOiDUQtfg1G58kN2Vfy5sjvROUzG0iB
hNnY8/j3C0uT/jRjUVGvK8Yp9iuxOARAgpdOEuPY5w7cEGRwSB+Hkk23mXK+m720bgk+rdF1Uh4V
eY8c/i6DpkayrdDEvj9pH3LqOfvD8cvCOem8qUcUvWnZxhjvVngTvUJcrqQnGnjTa7L5oHkFgeKN
ZTzYS2nUK1+5P07jGK+O0Ib6XjDNacPCc2UsLyo3KzJ7XY9g4y1i8lAbYGrw45plVtWrlZfxxPyR
cZWNCuBn5b3GdJ/AE0ON7sos7xjWkFoTBWHIixXKJrHY8jm3LR+woB3hNyL8KiY2O82JQw45cw82
Ry642PuK+U7tml4P5G9cHADXBMG+GgIxAkIZVOjYQyeZw++YQrdCEjTOHLR7QD2OH0gXblZl1oZg
I9/TQzmv+9ODkBhUYSb/7Lr39fCLrx9QJ2pU+jOaq0VRDAJ2MQfqGIeEVg2gVNBYzn3OXdOsyfTh
2P8iK/yAJdtvQ/Ri8DuxkHVkhZ4YrRLeFjIu745Fz/SXkeK8EE5k12gfqp7f6K/a9Low8IOzLF9x
6VYUWaprliY4T5TaNlRb8nbWIbwOORM9WhdWVGvDNRZx9XDRnETsT/KH9WoaIMBNUzCb/7CVMxuS
MuyDuYDk9s3f7BSWQ2peM8zB12xULdxQ9uWHIVMxRzzsduF3ofVD19AeEOV2BMxrgtaCiPTYcH1v
1o94hunKHFV9RT81zvJ+jTOtcHADtgO2syB0bfoAptysdf9hgeQs1EPWzve0kvax2sFFM8OOGaMi
OGg+WpY47gBNpVQYY2tFZOYXbg6QUEEQP7oGrfmkpMdEYabxbZ/swYuoxHjK2YK5NsqQ87VFc0ML
k5/S+dLhuGG+PIdNV5LTs2lZXcCSQ5TcEQcEYT9L+dsReuHNlbaKyh67lbJQGgyWslJqryepvlCS
aTZ5eIqrtTVG7oK4B+/DIA7WJ6Di+Qd7ClYXi0Ml9u8lZ3X/lOm5ibDzDPWA7squyBY8u1xcBNVU
J+ERoL0+P5AzM5WFXKxXQ0JRjoXWARLsr9mzKtRQkMif0e7TgrydwnyW7EwyM7/UpVSfVxf67kNP
pL45lbKUfqh/cCgxeeXgcMN//+Zm6BLlRZycbBj4zBGenx3v+cQVJOoyhreolHeeEUL9kwl5eopa
A5Wyq9/nSrDgXSxjk/O6nrNyU6WTP+2hN8dCXdOfld2mvMWWLynFrATLUYOn9VREi3Zur9iKHkEG
WJLpz7YmJ6OvmOZCSFkyBBaDm3LRGGyUrD8oQHvJCTemcTboBUTE+Muvo8wqCZLmXOZNPUmxnpf+
14uD/4/iUu4pMAL1o1Bt/wWJ5W02fijYRPGUHm4QBNrg1dlxgsuDgVL0GDexhkr48GiZQA+tNm5s
Y+WEv9GWHLix/LGPxoddCXJrRCS/1IjJgwEWkIM8/Pk45rJ2YJKJAfdJgdF3+2MgeKoW71GAWVwh
2lBqVeyouVH5QWJJSkWwMKNBDRpLf9IviQlQLOgK+c9lZmc0vzxrwWAqnAM+waEwmp7ecF4aal4T
D2XZyTm/HMUY4D44k/AVQh6WCOp3cdhPJ6CZx8U5yIa4VOUSJPu8TTQWwz63HLmuVGKmlgI9bJ9N
7+bwrw42j4EaPLJWv2gUk4gRa14uxFh8yDD8v8jeAglqmA8cioJdmnMzSdHSZZeEDAh5DrpraBrk
OaO54T9iTwS3Fqs5HM5D+NQMe5NwrgICC5hNU0BO+d7/0Q0evATm7L/DLn6RGypTprDMrgok7U8E
ZemfPHr4kI3MHwHbU0J6ANdhhdQAH7CmDNxzYuwm5iOFdXyqCzEwFamBDbAJN47cvBkKWoXRYdQJ
itioC2E2fPrQP3m4l7pqZ+0wA8bpGzVHbqJpC6UwqMFfJdUa+rVEoh//25ZtJAo9otnsZbpSyKG6
8RMF1tukzcmTAuHlEd3uaUhLbapLL19uAZ3OP8kudrSS67ZV2/EyijRFIo/CfjvfvrHoaTvMycT4
97zjf0YUybUqsFTNNI+YviHBfa/wxFVQTD0hWmGWOYKySCtLEBdCkXYAMZWLXLFz66AV4AMm2V2n
GsKlXiF8K3W4RfWzhIAydL6qy7KVD9Xe0Wrkv980RobdL+WhAgeoObPPrsJQcX60YJR1ciy5EKKo
pHMYuJSe3X4lkjAR4HElCcP2dqUkFSlb8GqjsFKLmpwAIIPDBZWgeRVQYWfp17FKq25o9GRYcBhi
E6zYLfqHckwGZ5a17MrygcMEzHQK1ysQNB+/x5ozuNTvXdn/p1HIHHCPQQDVkxk2tnh/R+nkXtaY
JIrLrWf15KNNcbvQUS5rsIZF4AJKyhttdzmmDVvNtiYS/AR8XTKgFHmwYBK5V04GPnnq+Y8VYb1T
dYFax+k2ghsZzbi1YZMq90QwpKCGyyfcPP1VCTQZV7fYrCxdJBBznNNAqHW+YgIDVkpHN9NFbs8F
qMY5FcRv4Ouv9xESHjXgh0PdLpLv839GRJ7S+nbLTQig948UWDX5Ucq6fuSbhd7C0RZVpmAIYPzz
agyF2CTtZBJ4FdxxCKw4dWV2y54JuJd962Ng5CF3Qnwfss3afVE5+UlS76S5VwIVt1eejyfy6OQW
f6hohegCTiypefmJOCfUhGGcsogn5rpmGUqRlOoh/HbYsDt/nrt+h/cAK1lwRfHtfIJAwvaIZQtg
tPDmJWFphrV5oUN0W3JFI0KuNTiyDWCk6IeOzsdRhzyIYF74VBQtoUctVY+zm6Exv78ss+trs9U9
UJwn6U8jiGN2sSj7YmxakrSwgBV6ksqhB2iuw2XUMrKLC5juAnvZmPLb0GSl1Jd078ik4VbXvG8y
IPCl8EPT2TR9a5zOzC4jyWjgRMIgy77WOrW3jfY9mYDwwjudEWZ9qGkOICUT+1WpGhhxdlxBpcVZ
ymvouipIJPrI8t49tBoDjtI6BSSHJWjabBuhzgXupZirpfUf0q1bEUH4p8GFBoqLcxLRUDsLz7B1
DZxY6DdWuwN4hdYyH6wyXmOrM3r0ITYuDdYrKF4X3yYgGifi0OfvlutF6P+cVAyONXiAdIYA7qlI
b5Xdru2es8Ow79kBEhEwwWX4NJizPH9YTZkrvdQdXk02X1199vR+0yv5itbBgveEoL6PvKfXkiTL
wMkTSd0BAWRU4MBWBbRMM41fn+pIrPyRe64+hNxTYFgAuyFJtXyYsDJlYzSn5vGE1OEqcb+eiuA4
oL67s0arPX7AN4+GIAd6g5N/WoGNQWJFYvFF+8YTfCy3Kub/1cxJv6gkGARoGumfRN/xdW66rEZR
eef0yfSu+jePeAsBXvu/RzZmIxCFyXKddXlkVv9u1zdFHZ5KAa77T5tOCbCG6YYfIOCwqINo9HLO
Id1aSPMvR95lPrJjcJufX12nvhq9Fnr3vix8+nbUFmRO1kknhDXgJHulLNTkszSYMN4BooEpx4Zj
FEyEp7GXfQ1ipW37SNw2+EC/uc6YsRuJqbUnomLSfn0imSEa0lUe4/33cwBu/YeeGYbzAtmANogl
Z+eSUVTeHD80SUZIVDcnNIhJgMMWXVak4xpLqqtjEA5Fuxt0T04H9V9f9zJbHX7X101Dk+QSwsir
kBf+rwQm/dqzeS3afEJSfwRm5jh7lpgehE7LfHX3K6cO6NTQqJ5rPD4el9N4LaJKh1bIr2FsW4zq
waDJsm9zVNM20nQVnuLxhJs5PqcGfYxzM9Qr3FBu6stxUf13zW3nND8Eb4k96a+KbY0cckFvk+ws
rrVskpswrTTA+69izvDjnoMC2NKfUcTG/xpLtl+zhWVApCtOxJaU0TsSgZdTx0JOdwI8ENufJ+a9
ApnhR2wX6b/8TEPRGUVPUypJ8r5IOgKvr8jukZhbxrUqNWAM4fjVjUq0YKLQqfaNNB3cO7gi4N2c
NxHUHKMZPsAD6XBJiW7oyrl5rWuq9k9F+5qREdeu8iGpakDKd0wD+YLavI1bhLYqFpGda7SVG1xM
x218rdgPDPBz3/kL50HzU1c3sGD1Hsvi+G26QQ+wowgGBnlx3szpiw9klR/6i0qeBbny7DmNUtnE
LqsFWsvEn2RPVn2/n4GVGQqaPXMH4BYLkBEUXCXEXhfvZkaIwbNAcyc5wOFzX+dr2EMPh/p+Fe2U
xGHB2XbHXtfBMhjaut+hRcGUGd96F6eCi17+zC9ZEoX1AeXJYJoQR5gvg/MNt5XfUoMOeK/ZZufw
+hP9gPSW/6s/hQ31pfuq4jbm3pBW8Ah0wvli+pdrmUbqmxoS6HGDAqvMnVoaJ6SqTs4JeIsZHnvT
OpN4z32NrBjQ+jpjPp/r2HeEmO11vGakgHL/fwluW19lEkJYfDYRhooLGafeUQtqTHPCuNOuAvJ/
KhqbX4lgM0oGyH6wcvg+Fs9pstoB4X5IRMNLfAPtnRk0ggWit9ZmGW6obAxGZHXW/hYehCDW42CP
v+kpOJs3P28eNXhz0MM/IIxA0fXX/NjitZUMNpOFfefeIxSwJEZg6ADWX8NwGhtw0BZQ9YUZjvX8
TMOBvXuJYDPoFQ2utdBZZl3qUZV6unaOE3I67AN6T0imA7/Aveu4FAtcV7XcKQrc6JtH38k3e7EV
TFVckbc+J6M93oe/wimTWpW5vVMB+p2JHdSV0P3gZ6gmH/H57BDEMYAnXSy5PEyn9XgkB2auACwz
eWf45WvrY+hrAEvfa/hrgQypKchauwTXg8m2rBSxDJUBMk7q4s5ryg6yAgWNrm4+bY/81QSy017E
OaA2Gz/WN89kHkOfvtriJiA1pX7X/fYtZmZeOcc1WpQ/kT64Ys2dJfAtrF8H0GdGMa+Ae8oyc5se
6MAs2/+4QY2D0Zw0/AtxB2UfR2QCiie9O1sJ2ygtA3pukeuxVetXFhkHa6V+DN4jxBHnli1j3AB9
/LDQBt82D5+nYhh/eRfrOiJ6cFqDynIOybhm4pd9xrI7mK8gqR1FcSiMgQ9tlYp+v7M7E7vbq6l7
bQTa8e3dNVF/VenxOtBHAE7qkTFm/GBTl91O2FRINplswqXCyldsSleZ85U8/Hq13ogY+VAAqZza
jH+ru0DSTZSSJwLqyocvFgcgQp4SsgJd0+enBtjQbFsKObEw0vrb6RNIV8KfJColorHCOG6O3X9N
SSUS+FGNQFf65TJP4arnTwwSDPB9tR8EexHcYEH0ihWjJk33YrEM9kS2rArlv/KzWFYu4qM1Vsx5
wLbif57FY+t/GsYOM1E4OyZbeBldJWmArtpkXSah/OVl1wiaQi6LFavF/sXw2zTUGH4R/SOQvDD/
aooy1i+2WLNs8Q4meQ0Qj32QUsAUdsF5mxehD5sGdplf7CTvRAmao7irvc7/pv+Z22R+4UOH97/9
VE1vSL8FH/6CRX2ILqepet9uwoKj3eH5CS92VUiqY+cVS/MLqVuzhHmAXZE8dKMvLJBsbiqpR0OY
LBgjsDx+eWhnOdCnSNNohv8aUR+rNMHHCzh/DYPrWV1y2ev+2D4Ul2u8Ym3dDBNQKLwGjzUDBwHW
LfzI3MTrglpGQKbazMU7sIMI3I/5r48qLLgFX2/aBPi1U3IC0FMkZTKXEyd4eEciYlATV1QEd+eO
X84g+LWSAZhS2J7hz6e5cWWpJt+YqcG8dk77+dLHnQPCZibbLvbalVrltnYv1HXFrbsr+203euOs
lKr1z7/aOxsPW3WJk8g3d29xlDH/GHEm77SGFEmsuCmSL42aZpsazPkhPT7gyiM2UIOZYfpY6G1H
VTE7z+tz+g6AbUpWyMnAA420A1Xi9fWLsN5Vp32UlwaSb/imLNZPFJr8vE/nr612/33ihDTx5pgQ
HZ3j69T41Bx5RZup2rYYnL2DzdWP5MfvjPU/yEyM+1dZrT7AZRfcXze7SbqkDzrP7Y4Bwom6Y7u7
hGB6DW52Tm3jV9cSsg7M+kHCoRVt2Vm4xT7aJwZM/4KjiBCyjNiWY4DO1YM+PlLp0cyFGLtbGJms
wpqOy7+FUrZOkwJI/YObbdlUx6p0IfbfMIwW0ZU7yGU9EeQ202NAz3egEY/gu+9uojIe4A/XiUUl
p1JwwDjVVFDwYQ39TNdNDvj6bsR4fEOWyqfiMGEjFb991MPS5DbAVgJSipt0WAP1n/BlmhXByYBq
MoeIymD+TvKBvexL4U5C+AqJ1GBPwou7bi7SW3W3EVpfaj2E1gKMWS9vwcPK+BErFvbIhttRq0fj
7DFcjxqPrEwXeEAKgaDyn1tED7XwmgQxah6dIsEvlmis6kjNOcFGofkwpEceHUxxSeFJm8T3NjCr
Gsu5v+yOXPWogPECddq2Jr4mkjd79MASqtczbchyCdy4E6XJOZsnK5jmrbwB4ZJyguxNThuUoZbw
Xj8XnHEYLqg6D8zqv80yLiofwj43ynAGCXyv9kvTJyRpNhcVsjZryCuq+vxohE4MQSNUYb80ZZKL
Ii902BgQOVBwRGI3mv5Y8biXk4Al+Lumg0TuyVzZDkS14CtutOOzyKQ0nCFYhIgAyp+ul1t34fGw
tlGYotFIwtDzPCUd/WC4MX8x6cZkwtuLhowHuV66SaFX4W2mpeq8bRyTkuwqakYsAPyZ76asjjJk
qVE793H4W9glLYE0yFkmiw7xKVi70HS3c2AkAwzTjo0R5EHzVYjYDHp2uUmOXbT6/uDqDrXWNfLz
qYVuZf9Rzhz5ZhewNA/yocM2lCEy4MSnHujSMGHTw4IboRgs9buOETDpFgSdVw7vJ/Edr9Cuh/un
5aSETT8Nrbo1FerwaPg9gvSe4GY74d9/vWtcAwLJJfc8G5k+eB0LGEy3kcPwFFrfwqQZCkPa+/Qf
GpKXcvW5nTdh9reH8N/ypr3hbHMGKJgWfjNcoyU0JzPdOJ6KCUy7Rt/olIg1z3mFVENGVAzY1dZU
M/BL7ZAcAeTwcNn9wOrhNB0N61/hf/p0TWJU/oqTFbhZUxrSpu6E2pA7e5YFRvc5U10dVGcsw34E
+5kiwEIZ1pvgOMt+mg4z23Ami0mHHcSFocE3s6G4lE91E0TJwfhCwPXDYcQ3s5eV313VTzHmEChJ
agJBz9Ic1mXn8z4n5mU04xdegwAmaqJwYzhVAfc8/o0DFqXkoeCykgsX3U/Vk6upys29j6rtqj3G
cXYHIcngHA8ucc897FUkp69KvnpYyY6HM7lrFByY3BtvJm3KLYkOApI6FzI98DNDqfhTHmg07s3F
Te31jZyHIOGzCZAFAvVM9GtvE3u6QjxA/ipet/uKfhj74hrt4vtyjeMNLbv3kd5XlY/RpBktQOFK
+SPywVRcoUEiQcume0/gpIh9ub2iMudR6PYRXOseicyxucVmjgpOlHnNM4tQTQujRe44OtjLgaPb
xYPZMfyf1jvV6PLqzZd1zFWwv6Z4RCriau1ihevZeL6SeojXdz3+nn94WnQSBRkC8fyLmSIUDQwx
rVJeqivWwfIqMzFDlWbAFBqIzLHchYUtA4bTjiWDTGyb4NKmotWFGkg4/8/+neCb0M7LkR2Rk4VI
wigRMJu4MN4fvz4+mdMZ+xFM+Oxg5Qvj4BNx8+Xg7/3WCAmmYdJNIGHF0O5/qB5ra0BiTTDqtj3v
c9Fc6RuVsIb2Kul2HjdPMvXuKV1RmDu+iVMifsaidbmFsggf3AFoypY3qBaWTE4EDET56LJ4n82c
RzZKMgOdIu6Bk3digekwzBmakDfvuSDIOn6yHU/9v4ucc6GJSG8f0w9rg2dCMRvodilYxZ/+LAMg
iQKFyzYM9MKLMt8EcHfC2JJd8JGURsfPi3ZyPPvXTuoc2dXV/RleXIUjzqg9zEcJd+U8V0lV0XeT
rhia2Px67A2xWBjwRU4uAycZ2qvBeonFbWUiBE89HBRNELCuVUk9aD4gTmbrceYFxuwxgT9RlXpc
lwtG4ChLF4Sg0HQdZeFpb13ZE44mHzR+lbAlAW2C/icPC4DTlo75WCpfZ4lOGLU9YDkKwZwYC9+z
pua5BE6OVT0zwV36blD/XyR/fGGTXMMPHh2y11phXwbwdWgVVjxCFmUPyIQ0gKc+XCv40Bg0+zH6
DMqLMdjsKKlBZ3A+IpLcE1RYbihtefLgAtFIAn0QbMBL6p0aLH7kL7hp92O2rvMaUSHAauh03P88
VMdfAE5KG0SIfHiNyjCoeeT2UCSVr7HvITkKGH4r+Ow5qxJ/srCAqNSCGF8fbZ28jJ6tfTsGaNHF
Y/S2Vfy0HMWEAG+kI2o/5feM6BeP2ZUKHYbbuj1oscIZOeFAdGpIsGoqjVCKfVgmcn92o+v4/4/g
q4y8fFbvYE5/SsU8JzKN7s9LyV7FH0syKLRP05edoKXX/1A3SfOgLrgUtAvu0dPUcmh45+hkmtrx
WM6Xx6kwzVkZcADVNgS+oTG6YSLvnY8Vt7vXnQslEsEEzAgBHlVJqgGs/jDY4k0QUV1SLL6qAnxq
7Wng41YRz332dgXiOMNT3lcx23VZaRuPBfmdrKzRcieZOHDrrtIca+2uxruxEGRoADtOnSnIUgF6
Zp0wZ7OjBwAliqpEEd2uDw5Bn5V0xi2hf3pnlIN7TOXbg4Ub1+2dEJLnGJWpBU/R9B4VbNB7Syzf
q58NzgAowMunN+O7EGk9UFgmrd30CC3BNAfyMZv3JKhnN9ZPbsHF7LW0Ew7XCVQHyEjkqlPEG4jk
+npfX/ucv7pED4cLuf/yHcB1cTPMHsbDeh6nikJs8g/HHh2A7X4HugnsjTJ49ePVG6sJ4xoEQQeT
QAzYMB7hOXu6uHZ2c5qD4WWKSWirgKE+It5syw5gsxUc9NqAqqy6dvD8/uB7DZ+roid17CgVpksn
IlpwgC6BGOD27zpSFi7JiJRM36hhMUk+6Ln3jP4VKL9jSIGpEkjWp9zbbeSGCmSRhUeEbQpN/dyl
j0h3IW8uwTtyy9zAAMJxcwCpz+kKr4Sxocqea/iuxy+uhcECmY/UuHNuvRa8r+dCuca/fWdsP1mL
iAjUUokxCR4znuGLmCWj4JaADtr61aLOuQbOWvxw+vYJtyRrK2Gnl5bd6sgM7ViqOGXWP0WUkupt
kayeb5z0wxn0XHeeFNjNsSLmxTrAjhKYcP4/pvtdcsr5LbK4daUk+nQnOcbFNNHIdocux+8xeBZD
2E9TCNbrw+QTwakm0Gam7zdha4fXkcAASzrHfbUh0MqRMMiWGWsTDFLnlTYIIUo75gsC5OQm+iWQ
gaCnz/6IfxWmq6nriJwrWh3ELvznGMHuIvVZhrjczT1CDBCCz7IB4X+8SaLXX0f+D+3jSH8PcnRx
6xUeKE/biSUxxjUZYa0QuLy4xwyKsQJbyqcTfim1uyAH/A8f0nGa1MyCfHaQbQpAu0Phg57iMJIt
f738AMYUMpVsVuLaXFEMClOfvGQ41yjv8O9p0414VJJGIjPpqqV54zB0TbXfrAZVZwpliZ9UeZ+L
VJwqEDPnYOxfzPu2lCqkBUc1HbzSuclMllv7kau4dJ3B6FIq+Y1poPIZhuRerCRd4ZbwkbeGBp8q
s5mE5ZDT+xehh2d0UcysSxHV3et4LCIq7CDoI6ORUe3pPwhn17sc6NFlg7/zootVrU6ii//ulRHu
gLgHfFlWoVZgDgzc566dYqht4fjADewGRC6Srhhtbw4tRwjiMl8Vu4HZXA44808bWKG5vsGSWB4o
qGmVgao6mhtPvXcJOSR+qj5HrRJlPojlIOYtbAR1ATmHu3+c++i3AIfkGvllM2jYW3rvNq4i/zPR
Ghk2BJvrRTqcw8dj4FMaL5hljLeNCsm2BDzVHpCRRwOf9WnJDFJqU2yNNX85uw/p/WDkDGfTY9y9
/CCvf3UjjUYr3bVVNTlnge3wcyUac7Ys51NeUj12vDuATSdzc3M8X12K2nLs+XXCqc24CgBU4JAc
E5fR9E4EEGjhQ/9vJNzD9qnBAqZ24bruRTT3j7MEjjMPLaVdFZxRqhagv+BbdhtCH/HyR82NgAf0
G2vIZOaqIhE4rBQSCEqWnhAPQ+0YI+KPupf04svw0VyQbMOzLZ6ee6gITW3oEV2anOzL/iZToC8f
xEoDsLLmdaB6mTtWigzMMAsbnFHD1zlvAuxNpbgSqxd2Gy9p6IP3DUKE6DehkokLDKdzFTaHDqtE
cfx826zC5RF7X2Dk7Oekv7eh17teQ6QVQcXq28TDuElmFA9OEH2YiPAu6T8LgsSSL923el8BUucU
GoOGe09Gl5cMFduGmR8xs0cHcsUHx5heoVnQVGggSIFNMWtWctxhpJLLkSVDIx0QDRLDuvswCiex
8v/XNQ93TcUDE1PiG/miy4kiHOduatm+1HLqbFzSCVAQrXkjlMqab4XnSfgD51gA2nqE8N09LUry
z98v+k4DBZaoi21hMm0Ojuxg9CVFYW9Qh4OnJFVb3mP9J1469NnOnSrDDYfgyRCP5e/RSRj3YxnM
2SnQVmWsT9HXErAyTJ/b0eadTNTVoNG8WIOPvWGGUNYef+VFZw35p9+f1Hh2VLLYNP45KIx7+g1T
2ubZdyZJthnwG7ynVk4WkmX46vBgoKxST71rjVX4wkF4ZAgxNFK9TSgvNw5HSVmE+ENBw4d64Jyk
Qc9w5crEKImjhu0eOb+s2YU9JivrPcKdt/N+X8LHcVazZAXUhvgpuWKTbndL///mjB+MljJyhO3N
4LK6GqTgFFtWgTgc2n+IUQ6qMXMOEbU+llaH7wtapBoklp5CQeUkDu1zkyFXl1clP240V3/kcHl3
mvB8oeth0bzPZ93GsdlHdGrYeB2uY8I6UNi1JRt3YwYO0QKbwUkBturO3WflkxOSc2bd4BrpTi3E
fNbZLqi8KkeJAXGfjTRsv3zPoTzLs1lIwPvzl0q2Nu0OOAWgBHZEujKLd/uLKJ0wW9pc+m60IkFX
lSLXn58udJmbMVGFwI6+pc31jtomggGA03pt6TXVdJMOad1m+hK9KUNirhXnphVVVx6anFVOU/cT
uQbtWGWzz94FYeNyDn3kmWWPPzeMqJ99RAZGRUDEmAx+qfvOwAUBLjOW3GPVLdGbZbtarYFtJKAf
A4vxXExoa/5skkK9HTBA9R330lewRobWz3aJkwJppYOuU6z77+ksuNVFpcgr3zlRp4CwiPpL5oTe
vTvZ5UAwPbJzLewd7rhTuYa2JmdR8wlngJOmKCtEl3ZDiSsv3waAtW4e12lxUWwTPGFuhhkRKrmb
CDuAfzCe8idUkRuRdUjdsVBNeTxKWJBWQi42XawqeCJlzFgUG6DUKuuz+OtyqFhA6TQU3PWqyxI+
z9jtvVRPEqydwmRQE24vK3r/AuYmwLErsZrlw/DpqwSKEPZchXCK/koTWjGm7gHtmpkqrqngrNs6
iN9RKbhp2jHJ++eC4I4cL6y/f8pdxLJb2CV/SWAuIfXjghAAqvTmQT82HCWEAs8+g2eWkzsHHoeb
b0tPjYNn93mGWz9eJHEnIsZkLQuvxVqA8agoy/Mij2JPp2a5ToDr/A9CualgL/cnJy/Dxw5xRQ3e
vEIS4AvvZ2E5yVKCSBFwalOiNjuJPt/jX/M/Ts6m56EIuLi/ApamzjMVEB7O1z1f/QXarNAL0t2I
qIjrQK4/E9gU11/zLT+lv8oEypFAwUe24zX4T9tYCuzqoZKHwxk3ePcMOE9/FGWwi4tkK6jzL8iT
1CufeMwUoGnTsrVzntyVlxEADQRxsSonUjLlpKmDyZf7l8Ra8Xk7bqFs/1jZSzQpqXQ0tWdhzbra
IShQAd8S0NO3CNdDs0uiehGp+zSRTy2zguogNUbRjtk0YFhVUmAxpF371V+Bu8M0PYZjbuoiyD9S
4xtrCXIBavwchz/udmu4zm30jIOc8qMsa/3cKx+KuCB2rJ82Gg7KZ8wT8hAmTwnbp8DebykXUB9N
rLFlnpjcFIRzDKLgtpxlqmx6ZJS6cZUlhg/dpv5DCDvMxc3VKGTxkWIrXmJO4chbXtuJVmMJUv/6
mYcDBJVPV556RGPPcXdbrkb+fJRtjsQHsFMhrn1ld/9ljJYobpT1roYVvzMulsRBuIGwBb8qonDM
7ZeoB0sDr6QD/vOt9qSPuEu4HzkxHjy6j+HQ1SJ0/R85cdxcQOfDAdjvBNJ97v3ax9pxLLDdemk4
APJHgy5Jfx+SpVRDF8ZtUeyZTr+QiIDzkZEgrNL9FzRH2lvMV/Q6aLAlxcLPyswlRf+To5vgxqc9
lpbCmOeETTXaXJes6RbZw36bupTRDbm5Bxc8P45de+qXGmaLuup37e/TUBM5wKFQRXEPMBKNgwZ4
IhvlqX7p5ZOAu+bE6Cr4qHd2XrJ0mNYjehMahXm4taP9IgxJRTl/XoP+MIoUb6vyMQMPU0QoKWMh
ruuIPrizyX4aUkZUgQoAk/Unl/IgK23bjfr0Q1uzeIEgsQiYakwVdet7Oyuzqztj2VN9n73reS4K
awn3NYBBdQhlhVQkLgAJXtjJBDxHeBDO4NxvXy1rPSmHNSmP4rkPbqr0sWuehqeNrvyLgGpaF/E8
2o8ep81h7rkPUGCweyGd0GuR/b7TEk5QyLtMDWclATnmOWfFh39dBJnSm2C/0cb7bhWEltdOkwf9
Ki3GNhMCzY3qCCcegjKJzZuCtGenVQt6GE/2FV7po0LDeim/nI1vH7EiKoqAHZzuH/ToWdiMb243
WFPcLQPRnGUc0oX15yhLtbXYA/bK9p+yOTybyx/4+9Ei+uPoHNxwOttCiUHkHHPLb+YE1OVcIqNf
CKbBYykmn5+0cilsxDS5fLyLhh2qD/OxQeAV4xYwlk7v5PNHNmqg2mwcvhtqzgQyUpVRXs3HTA9u
I9+QDcOhlxuGVxHlKzNR6SgvVukY+KcwZK1xAs7fhdROBL1m1TngQ9TrGHowaZawgibMew+Nr/H1
v/41Qq1/wz2hUTVy31Cc7/81JOUEWb6VQmKxwUSOdmRQ5s1Ee3cDyDwL3cohkrT8Mr3tueS243cL
/J1++SfcuY0Q9FzPG+FrfLH0m+DYrO2cqmfz4S6O1AGa+2tbEv9vLwARSPwzlZw4d2ydYfxLKLj8
O5CrIsXWHoaB9r6X45dXj9D+kg4/blN+mr4ZJ6Wg7EapLv53RBtwlFrRrqJ2FUhuFta+Qqb3udfx
M11SPGYMsMhCFUyWGfddIbMQLnqxOYxwdbh+4JXLH0WxIYPSPg8ujfHLMvdpx8k/r6fLMnJ4G2PS
y6YhdOE8X6MGI9XlOpwj1FQoC7NFe0+FSdu8sBH2LAnZ2FSyRi2APzTdSFqLxL5GVDeH24QkW3J5
U7OskR4VumQYhZgeLW6pe5zITY3FZXsXkpWh3mR1QO1CY8Tn2hTkxCaFs0p/RPLwBO6LDNrMgzTd
VvwCb4deAS3MTHfDSJBNiVOsvIADMP0YrMLWyU9CCcw7T9C3+oi4zJQGl9kzqI/n4ZhfniKNuQxQ
bDFmdMBe+EzAN32Ft+56jqii/MbPYrW62XtQK195hZfIVSHIKr160yHQzACcUCwFCKk04puIRgfS
F+HrySiB1bBBl4UU1Ocgyky5KC0GoGU41TcK3WoLZmdxRh9FeG5G8Bm1YjF60MfA063GZn5yMXpb
VW0By5vO4ecOZfY2mgb1yYPFYtfsACo9Ls1+HlZ0N49v13bPek42UfMKaMPHqR9hnPsv5V/i19dy
/Qemnjp+O5VTDOAxYF3gFf80WkiCptwOj2dMFV+Z8b0h041Vw/7JZ7T3XEphpTEXE4fVd/IbjLvX
KzLwhG6aPjkz53V6ygnTivQ8Cz8pP7Q1C7/iFe1XvYWRlpsN7FyEbiHJ1e4zaAoyMVJSEPc21mYy
pP0ZcVty5ZGG4U7/0HIqAzS4LDvb4HFlRyPyv+fRF5epbVuJNfXitnlv3GZ+AOyUluZkwSGFQaFD
T+9WsAqRJmDnndpY7Y9hfX6oTiip0h6f5xoEqX/vcvpf3tMHWnroX0yTWECnZuP4mYkoKA4VzhtP
0tu8QQUvyQKJhgXoYQgCyqI6atiRjnhywntURlhkU8X/IN9G/68CvR3AGFFb2o09qUeSO/ZVZ/dz
vUq58lV2h21AvPWCt29M6UjJJehLLDr3Vb1bTF1h7vgxlKR/eR/Zf+hZO3kAcRUGTTPRik4mMmfm
NF9V3oXnKCgRuVJ1akTt3TiVn+6ySmhgEUt2fIqCPrOpDJfByY4eelTOIV/2lu37PJlJ7eGZsaPg
wjrm3CnDdjXTTP4gEaJqv0ZXYdli4muiVTmXBdBDBdovzMHArhwC2n3oYUVkXb7t3Wk8X1EGmZz0
Iq8fOo5WG3BJdFD4t0N7TNuKHFDRFueB45Vsle8YJeUhJ5BB5xlRoEOwF/Ajw8X5qJUOTMsXLYR3
aH7YvY3D43UUQzl5WVUzr+FBPwMB0JDDcaSOg9QtqKusxA0sbjLwfS+CoY04oOlDnvkESiq4/ADR
X4V863TiBBP4B2i4BWk858pAi7NHqv/SiXpbfShV/H2BvDnpOi+Cvt0stdCqCNUSx09+RnqZz0NS
s1vZDBqUFErzaQdwmGRWRvabCJQMFBS+Ot2C4MRe+F5OlpN/Vz2btMt7atkmNeEA8Sq8FX8vk9qe
u5fbyRe8DHnYqIz2oH/EyAUZG4LX2REgdqZkN4tM1x51otiFrWUAJuVld2XGpNIP72XgdH/2nPbJ
9YuubWD4I9Jt4myIiNgiiw+3gdDvkmlFm4Kq/CkpEmXuzB67Z7DjjSfUnWc1HPc2/uZIz2W6U4WX
NbPhnk1qr/jZH1qnkv509GJlXDsjC5sxMLhI8tnpcXGWf6XdmYOCIvE5YlzmWaZSQaMjBhYHP7Q7
5oz07qtzLpkyza9eX7cUSKinc+ugFnXQ+QMyav5j7MV8RMiONodMJj5L/N6Gg89nJSbmNciNK8UI
pwasgPeDFzynzx/hj2paNLd1WemHRgOPRz4B/tjNMd9UPV6fy9arMSYRl2BIrn4plxWyrg8e/pQp
ECUksEqeAjn+xj3WUJhDdTLHyGbRwNi8sr76patawXlFg38ZQFXAjeIK01XXRG7aaGJkM1AtFo4j
AarNTqyUOpKdMeEjFLAA0OwqEATV0aaAuxnBBP2kIBTuOrFnIW8Nx+ekAKUSHednHDl09YdYCD09
uXKXFHqBlb7vibsx3tfuHGOkw+zZDUctAOQfDCDo0YQPndbmyRJRRgR1Uat1LfIR6/onmv3bjue1
twTDeIVVwJV4NsNvZsayVPQiE1wVQwDbkHzjF6K5kacmHOYReMdJrYsxnU/aehna4a4yTk+t+UYU
T1vL3aUh/SwAEqilZtNq78/jjfYtjut+D0ewO5za35DeemTXQdGnn+xJn+ZsPQ5o4GXNrzVYLnwQ
/tjyCZ0uWyM7DuOA1FVvvvIHITuEo+ZMiM/6qa+ek8v2l1V/6Sghnb5QVhyRSt62uw0fgBe7Mm3a
xiKQ8Rzkwv9TagB8dWWkCsIULtJ2Pw3DSiae43cA+hlpUJvSt9W6DTYQemRucIEFbYK6Biqjt9vu
zb9w871BbziMnNCkIaPiNN5aM9j13ltcO/MQYyXuSH5WPw/j/j5e3zOCPTiLb2kZb+N2qjUF6a3V
v9pTE0z+je88mmKWZIxKn7KsGM3+Py8LeBPvR1/Mjs56l1nIpUeD91GpFth6/E/j2ruYyzRcFRIN
+C3ihzTRWX7HNeIqo+ZnfmR/qZnInV2MkAG3uiFx9jbQc7SYzczqwglF7uxq7sB90u5l5qLjN5pM
npgGIgsIoQUz9Z606nPvsqbvXCZlm22br5zqa7DvFpRs3aPe33I7W8Amb/jMgnGEy0qoncfbcyMN
KHlWgHWyby/pRvU76pIubbaPxXfEGvvygDN364JCUb/sSGtRAmp5FNb/abNwKvwRqgpRy0YCaUjL
/kSAsRqN6QWM96pXgZMy3Bj/9jt6nG37a8qSDKTOc3XgKgiteLP60jLuoM0ipYMXc8Mjg0CCka4M
W9CfMmZ7z1cKnegy/lpSAROZs5es5BqsgvPdo4vUvUwF9T5kLaLQrScqImOcSBilTe7P2sXk9Fup
MLmLxSSS6AeEtsBXgAPiNmjuX4yPEpVD/wTFC7h5Xq5qciQb1lpx3r91jQu2FXxFtaS4zoc3JWNX
vg6US2GbVkxWApU+875CzxMWyTrej9FbJYrhpkTcnnWpaqhvrgJk4FRzna1u1mP9rR7wM1qvvOiO
DMDGcW4/+6+QE+FLx5OeY/dJVV4vzSzSi7PNpWj9FSqUrmsyZgXYotAGIJVVjgswupdWyK7gwUuK
+O7UAoK/AySOGtvpxqZ0nxXdKVvC4Gvl3OH38oBbhLsWWLJUxzHMbxBJ24YDVQCguTL6eBiRwzTM
iNIBBXqy4FAtS0iVEpU3XCWS9/xx02B9Ojgbjl8w5aCkUjwjUHwhu1b0XEBWw2gl7y/Q2FUSgEh3
SV7BB78uhCMGhfQxoQpWQVOEi/7+r7w65Jwjp7+wWCj96Pi5zbCUOln7VeWg2rRXfS6g/MHeBHEs
3OC4YHXX5HLfNILIUHsmquB0oubsLuDiBaIHcsHr7OAW8Q9zy0z2xAuF3SRz0C0E+rjnwJRm4LsK
cO1Ypa0eH4JzHX6qqYR1nLq0idCgpQMgbdKb34v0efQXXvcnp4DIJLx5ekxYZ1XjGlwXGfW1VYAG
ioZ2FHQNP2OIOrGkEW7ChzyxdSc0WunsdcmP7fOCNTQqMsxDKzzBHfBZNVy4qkyTtc1o7TIAs/gB
fa8/Zh3OrcT+dbZg6pdkFWs7Ioo1NixVK0oWDKnDN2RYZcIWrQ35pF4LQ/Ag0MN2YoBWv8CTz0qJ
KiMOLm15zbUDc85MUTCKI9eQWJR1zTVaKVWrj+cvdnhhq85l022qkHluVaKORScNcN6bEdO3pweh
JNO0GwCjlLDJWnr7gAHJ1ChyH8He7JE6Dn863PdYNe34Qv+VMY8BPcWrWoJwnpu/d8f4L4XoEfR0
O0RlOaU1ouUutUuWQY/Wz63o0mhdtdSgNyARzmwh2kJ8QbJIJPyqbxL7393Azi5rriUuEFrcKFPF
4/nKvT+ohBXkUEJ2JkXtMVtTByQ/H/cq3fvEKmQpmQahxw97uZVORxUdhnYGL9ynwIdwRzQgdPsq
O2eDEGZxEDuiqyfcC0VYwsIEbz/DnAfCS0zAP031hzhkAkqKNAo4tXXA/9Di7m1dg8j2vaY0RDHr
NKJsgGt2iwOugL8ECJsutWD9Bd116bL4zeW+mElFTRxgQp2IDHVyNh/XFZxUz4ZefnGrcPluVyko
SOd/ZUL67ntHYinkkKsawITSRy+5Qs9gMVc5JQQ8iQmf71xeOLXipy6s50md1PDBEj9jvMEvHkf8
M5iimNcbdJkWAZtMlsI3ot1HsxnNafvNeCiWHjnBieDwJfsiHojM3KsP5KZ47iNUAfAcksulXt/k
oW8XKRAOXZ1sNrMSZ7ijZdEtPcdmXSyjcporged4tHI6z8mSpN89ExHsAj8adP1F1LGFWf1rCOHe
R22AA8aoHEKzVkUB8Dl2c9cMvQMLzAaCvjQhRPLlWE/4eFERBOJgKSouJVzbdPdP9dM2EkOGqdSW
2e5itCSWMwpA+AifarNMPtEymaZkiVZ04NJS4fT5XRfENT0XdbnPOFOosb2ZALz3+Oew7SnuisRE
D983BlyfEWo0LpvKeA6niHnI6hhZ6oV0mv31Hk3H+YF+H2jJLop6INv+odpBuDDwhSoyANtWhGAN
uHAlu1joZ8gyDxVtq7o3KyBDOrDhj4A/879AZUmh3LgUGqzQvokg4SU+Oxelp2zai4EBCeQv4Ixo
JTtC0nCNjGgFDL/+d2aq8CTFFQa28WwVfHc2ncS58oWWpb0aBwn7psCFRpF5N1PDIZDZMVj9YEtq
nG8FDhw5UJSpwaZfEIz4DVGooIAKFC6ReU1x7oibijIMsD7zk+wVNh5v4DnDwOBpJgHOI5tyNIgn
0QFF5KgsD3La/55DaFBTI8tXDgeZSGld6iZe0pNbZJYq/UAgKKKpV7nnYnqQpu2ARimDZA/2fXc7
8e7uRYhYqGQWNN0VI+5UqpZCcET1Y9eVLG087k4oljdGSsW5zUK67Z5xjopmdL7muAJCc8MTywZu
fuWIra8CqmvvCYlFRH5o5Ow0Bn7txO9fQDCVjGDdoRaBwUvsITrFEDImDfPYsUbVAgVoKqvL6EJc
dUbNfG98jql4/H226RiROnckpWK8lgPXk3JQQNK4xqcXJ8yPFYZAd6v1FWp2z5FTBgXjqcem80+f
W0jXb/QjoeRG9u1hE0eWhK6Uw+h/995+z9KmemHkugikD4i8ZgudXdnEG94wlVvBZ8GhLdf8DKej
c627be8EEI1VA6C/WpSpT/BeTX7RjIZj5dEodpVy+QWCg3XQENr1/2HcfebFg85t2fyNVf0ztSZN
7r0ytmMZi09ftT8jwTg+7wf5v7QReZcFJxTmBTLZFDVuDipC3JlGecxWWTyJMt950tRHz379H4PR
uBiLxkLsOWifGdrEABRnROsiT68LHBZJVnZVHVPxb+98wXEdh62vJD2N0/GjZ3z2D8xxO3RBvjgo
AAftiX6Uk8HRFasBJgpVt6Sp5YLte296M/O1jImc3KI2nkXKdup4Lbc7FEXNja8NTWbh/B2v50RZ
GoRd0ZCixgbZTBgMRYgsUkLyLo0qWyv3DDbIbRfllsKJLI1L9VePE01+3PlLq9aedyV1Fr0gIdod
0/0DKX7vreF/Ip1zVAfx6gGiU0eaPj3eTIHofZIDevj4JoTKHJ2lkX6VKIYav9KFgMz8U3YwUG5p
P8rv0W24hM48OgG8g0NncSqOmw16PQCMHV942aqc79//kQGLXdpWA0A4pdKP3xwtv4E8FuCWa3MW
UOYmZtCj4RP9YrNQjjkKgmFrsI2fXzx0FVV36TSPsdGjng8TNNEqB165MOzjhiXiepufNLUj1/kM
89iM7mpBct7grC3shLEf624EcOHWUbQWBF6Dpw0Zg08JHtKMwSCkD+2Ej89POp3+mFN+8tdF/5vJ
5wbU/4VyZy17YFO6WxrMnKuEZFjMn9wFmd8V8kULJFHNYdPnXr7pdSNIxgzHpyHIpMQKtjaP5vVP
KINEjk1ikdXqcXhS1sc2f84LFSuXVbaciywbXKE+NM66VMcjauMRoBDxbhHW08F8oO1849YFqihv
kzCTL1DWBSzqPX91msH4JlOxrXHsnw9sXhii8sMinHtd+4a1hnojpRQ+HAsk1yzj3kIXwND5GgXr
6QF00rr5Td9NFEQXNCpgKNwNGSm11wHZ0PyD961SRtQWyg60XMbEPf9Piv/1s+Douxhe6GCD9DCi
nnqD6ewg7DhBVkqUa8Ckt1cFAbvRZRhFhyccL50bwZTM9iVM6vM2DIktRIq/QEICbpyGjAR5o2MR
Ts+1bihzYgzoj5YhfkK5obJaJh/9pwxeKfYCr/sbwxPqErFzFPG6Ml6S0EyrOKckYORtae9vL9fu
vc/RGYuttfwoUDEOTnQa4kLMCRkWnUvy/MI55/HwT/BRsWe8YZD6LT1JlmwQbZ3EuNN2Zd1LUS9c
c+w8owVXJYGosIid88YVRgI24iZxWyJppkdQppzMfxFwjQ7HA9/J6QuvI+ODDx0BZYwx4mnfX/9m
1f9UptZBNer6+8k5Dir/+FskY8zdA2EKd0wAZy/H/boiJ5M6YzgiVHgnRZkndwd84brHgAqCdxYL
VjFMWxsWlc3lPsshK5qejrwLQbdcCuLlfElHOCT3x6KD5YUXLRu1E5yNekQjUNLb6K3Z+RxXKlBm
QVbfpqdDMELHJ5S+rSQX2Bs7yGqxsbghuoZWbulSDBPL2Fl7bUoTn754DgkhWWyRFy4fKJeJgtST
xcNg+yAPIvWx8+ijNlYOkZ9l3981yWY/ZLPHBZPXvbF/a0wGA4OVWhfXyEZsLz7bz3M4WXuIcY+/
gNNoDkV+1w8Nxt6ZWHZJfzqT5heocGH5yQuTteQvmWCQVmsiEqwEcAyR/PB0VeajyDZYRcQ1zqJU
hMWFSXfrveqoWC0Q8mjHHSjk7nXz+onRGiP7bjfzopZkhgK01RzlV/XYdHEi/Z8onkL18cDK1qHh
0gI1oOjlg1V3UmyWI5GDRKXKFcUHdqeFfsH6G/0PLLBkmcqQOjg+jlkRM7bFYDmLPczQ+QeNh7lC
6MmO8QKUOpDbnbnEYf4JCpkEV+FwSpTS4t7tDxfBjKzBNgCzB1rOVsbPZ/nP+KqlbIfVc5m5hrsE
MVu1zB3xXCTGjS7KR2YCu2hDs7VCe8TJrPJH/7BpVn3pcl5w6+QgZePwZC0I64IKagbEmgr5rXsU
4irzXwtbMaBAW26KEsn+y/y+FM1HNbmAy8oKuDMp041sgKAwZXrFn0xvtMm47K49rZnmj5CgaUbQ
wGjsTcqZ89xRwOJlwlzDYuhmQjHsAl9pC68fS+obPSq3/dndvxLuCeaB/1UJWhg0GT2HTYAu5oFa
uz3y56kjDZcYDMR1QTnzO0vnO6AlSK+LELjANXsR57jUwYlfyhNhzQoiR5vfEcAorr9M55RSlDmF
rKw/Y28grNqDOe3cKEnPH28/q3VvHnYoeCo4aMup/aBQav/njlyjDFS24cu2ij/cSpU9AvN5ouxi
/fDWMzsEaG6bJaNmTGaEIr9R4QwaBja4jff8pVbXVvtZtEKwHLuk0bYQaRNGGcn1UHxba5AKMd54
hyfoPH8g2rtd4wM+0OR6m43LL1oGQo2JoZ29Humqg5NkVYvnpFWTAmqoYyoushlWVZP7huRzpo0L
K9yU39BuqmxOXEmFP9ik8eeCleZCcIyXK5Ls1N3XAnTeRU4nycV2dlN8AZfC4rJiIUnR+pPDsnRu
rCuYnyFSrYDzNxTN2jOY9blOKdYviKgzxphEsMn7QZHgIMAt2oIIIzOGQaPmGUkiSC2DbR/J9yq4
ke9IGXspZrJhn/4ZDmpZM5Y4TFs3wta7JR76ZFl0EnhwUmSKo2gZzCVho5MFALuwXuB+KL1cgDse
kPvDraxpqP7rJkZ9WmLQ/rEqfXy9euaXcPsAimx2si1G4qns78xz719/tuPNTxhH7vEuHxYRZ6ay
/GWRlpG4b8ZRUr3+Nz4E6IV0QSoHqXZzrj+PN4PafpDn1egEbWo1GEQLO6TCrMZt6Yff5I9ZYVI9
19B9Kdr4HxiiDn6ghH36ewZG3UXiK3ibKePVlpfJE03k1V+Gv+x5F9kNyP3GAesV0Y1MXjY7+UJb
hgVM33w3Xe0pOhF7/LMVXf22QkAXqqoJbVvdu3DbMuRC5mHfOzeS878Hn6VRgTuPf1hy9gquvMcG
ZoqZFJU5GtT51MkBucU3LBQuqLPDpREFsY+yxouZDhxPUOf0H5ddX2g8xFAcVYAWLKvwZKc5EQTz
6oZA8se9tWJyGWW2nzXA9jroFgYPvddWl4cchZ5DfT6mwWt5utYgvv8PN8Zi43a2kaqoJoQVyCB9
kFDgMGGckP2yiP7TYqHTeOLMCPfcTug/954WMCl9HB8lTlx74Ef2x/jc3i1gxcnmMBZapTuHgxuv
Nlxa5TkilYI0O7ONT13tZXURXp8nenpxJCEWztQCIIZlR6nfNXrHPGw+c8Khbaq0zufmSvaXtN+X
veAh/lGDq11TuaF4NKwh3HUQVycSaMwrb4TxyS7vJBPRiWUzUdmFeG3zaIpBH5yCnwFnQKQjW75u
tEfLmsWamN96gkWIRd4nA+k/CQZrgc2Qn0Q86P74RN2JjwHSFQru1ypoAJaDyVRC6pfvP4YxG3Ka
YTMrGvLJvABOigi0wIdm3cBuCNIGvGWFo94GqbaddwUxdyR+Rn3GsMZ9vAD22acaLC6FkgzumEVW
BbQ+ZhcCTN8LLgyic5WEofHgYGJBlaTFpUCUUowX5uhlIp9/FRFvvGokui9OaXrvqpceCUElDwrU
r/RUTYmGSxISNMLTS7/9pzIULu4mbC7FEogAm4rBgnpkO80WJmFot8BIEdyr4hIAoMpQQQHyrfNX
/iEwaCU3NixAHEhhlx115K8tgi7mA2Oe7fPhKJ7edrpSJU3V5q/MzCcj5zqbbfQSzEcBAUtTCgJb
PIuChfW/5poldMzGSOdKatSe7T3ppIyn1zVrPLDIzLEaXWJaLF5okwg3bWDC6taTfbamXa3ckiJF
T8+iqfeU3T9t0Zt3ZQh0SkbNuyOq6piB9PvGtY3V4FC3eujUXGgAlkJxozc20fgp9/5YIp6HKCKW
Hcqy/brdtkYXWH1zE/AdvWpMRDJmSrMZEVf2kEaztk+1jZ3Y76lOw2ol1c5UZWw4/rR2OzBJlkQo
5tBiaoDrjBeoU3V27KKBpFcF3YVIUZyuKb1fB0K35281Vr8ncTofndIdoU6A5qqXC3UjdXfpb4Fp
gUUurcFddQb2RlAlDqAcopYvqzhurIsOr4NOYOa5Lzy3lDmEPN0WU/oIij3wI5rWu4O6gh7qVsgB
TvsMJky+zshJnq4w4HXsYaqdkfn3+X8RIKdB2S1Wnyjfvn0F6sCog0w2EOtD1cU0Afjr9glhKg/O
mwDGHeTYX+T0Q8lJg5rslgvK0TDGq4UrlThCGQ1rPEGBinMiMRPpTZTKgQJM92efGLeOKJodKAkG
hZB+jEbMmqkXIWGjA8brWfZnNy/RbRzZUavBspMyoNWqNGUfUasEkJ5W0mmVHYT+Pu7YMamF000c
pmKVPV6FwddMPc5bJ3ylhKGXI1KFCCjB0cc3py1urtkMMx3YL9fPBKhlQG86KkRjpaU97aOiW8ut
glAL61c/7VVRzsKHR2CUoyAx7dRn/ciWP+hL8ppZTPz1Odi6GHGRqMUbAyqge72nu2i9dl/PfLQC
MpAW9LJTXsrquai3SZrxDQnYGy+8SUJEdvNSFDXcQNjxnqrvMZr0neUffhmXrYV1C2x4X/5HVlWV
dlggglOYTV9Rfxcuo8KHLSXH+DrsiY1E41wGj09gidS+kyocgQn5TtkcG2MBNDmASXRLgtdRe52g
AprYAMb0YkDBU3eSeKVLvW4CKhkObETX8w1U8m7Dn7/t5pfAl/Qod1U/c0DohdfJcgpbr6akW8Kj
gIaRBmLkhVGRvZi4+w6lWve1mBhSSU1+n7WoZ0eujdpSfJbGtpls+smyOjKTQT5NprEvOXh0d20D
YCX6gollj8ySeMK9p//77MEfniM9rclNlQFfwGLBapnHbkNwUkaRNFupgNV9pxxgfjDyUzxHUhoP
OZDzUsCziwG/fLGoTvD6js5d+noFxpXaVrrYFFzfjXxmmlDwBRth5bUTmfaLLlKrjCHKV/8+I68x
RgCnK8ZENLT2II063doGQ6SxydJDd401j+FfGATKpLX7Y1jR5HrdrxfVCV37PAMUCPEm8OdbrSN+
tkmjl4Rimrw9nL7fSu92pEklB23rTPwAKCYfE9Gc7Q1VA3jso3xI9h5ZwDbEFtU9yjdf0zGTt8sK
UHLYO2Ljfo+4ldI9wIzN16kMBF2TJxVSUuW3bSWB+6zzXQbEbRnt63+UeddV/DJcJK0TX+6A80u9
KuLs0VD55u8bR+D/UrZtdHYFESJ7XEwboh8+HeaOxo5QtV4dkSdkhsBzvbJmBk8s1uNdzGPkQJKV
4bcWpEOeBbnXEvh4xWlOgiU1bgG9p6KSuO6as9nbOGVfIXfQd/Ghm5iWzwzdhgusbm75Zj1OOlTW
8vPi1+ZG5XK5YkzRb9bkqIKfUPs4+2s6v6sVeQPo06geMh3sDuC71sxplOCEBtsjjvj/0u2PEh84
sc1xmZmUZ4g1+YhDbTonFBqSyop+FgiMBdLdxdwBsvHFSXfOBaZaya6MEksdx1/XJvVyCPkL9sv+
fXYgM4jH3XDztoqe3iSGNwyyxk6b7LKim0sEO9vKGiNmzrbNptxxoHmTpPwEiKV2my2BOFBnAsmP
bc3Ivsix6HFpGxC5iTW3vGCHD9AEu5W8MPWtJz0CA9bsfb2OqEhLUVxxbugioWtj6ePugykqMahK
9Nat/3Kpkq+s0siIffebEky01grGdGkgSiW8TEOHqQQoouZw9X0evPHbmzjoPGeJjsNJCC5C4ImO
VHIm1wJP4kvLxH9FBGMC0s2e5huvD1lqO/wXo6aK5+ZAR2xv/f3gN8XkMTz7v6TvKQJ+8qhNaZBu
vnMfqaI8GGiaH/6+cJg7a2GluKMKAFGjoLqz9ImNxjJvzXWey5hg60+9ZVQyL6GrJsBP+V0YAstv
uz9MKjh5ezPT8IYC5ktZTo7znm6cpq0Hpx0Q/WgCqvfD+YbeRmcNIXg3sJy+6gOTY5DhRNl5i6Er
BRz54p0lXZVj1sMJI/MMMcHT7U/bkesoR6IRsPOfG0Tnj2vai6ysv1F4HDgJAGalDd62WTv0o+7W
vQTdtwlqS2u+jqVNG1UxteGktKc6Btflt7JXUo5JYjsfiyfHt46VIahyR397aq47L6nmKwmj6hTZ
f6AQfCoIWNSiT2TdtoTqBVuX2gld6Lg0mjeEeoEFTLdITKgrPLxr0LYlbcvJ9HvpEirWMDTV/zNf
zh2bRDdF+awNeojiYCAL/55VfPxDXMpB2ygAmbB06q/wmNLw3A9L5xfjYWhGFuBGIPZabVfpOQf1
qjGl2C/M++xSeuytSFHQ5OeB/Cw4NKyXDu8lO7iz3Co6DmjSm3FrTPM7oNXeR4HyvhT4vD4QDVs2
EMPvcv7NlramgOocIUNlaZdbpJPSDcf7UkE4bfDlfdJtfroGe+VwqG6Hcc/TIFqpAsCLq3h3y0si
huNiNLalrE7vjIzOl0uekNUM9VOLCkBRYBkDZIU0CtdeCtbZ7MtAxI4q1EJ6G/M4sMq8qNUGBfZ5
wcG2n86Beir62ObbWMfR4P9XesgWDDtnapWpwWb/GWubFS8kwqQs//vb6BD+H32FoK5zfwC0WrQW
KogRqTEPNFHpNqLPc367SJWHLHvFK3ign9ijlywKp34olHK+uyHgLurtqZbwNJTEUUfXw9EmtEYJ
+UrCjSYhIbgVJ/IDkaXbKMcDl9uRV9XG22BSXozg/T9/cxWxZmuutofQZ6BBhlICg1Ox5CrhG57e
wa9iZIPL0z/uPav2F11jcq3Ja+qzCr/vmM21Y7/0Wqn2FfJkVYP8zVdcBtAX2EIQ4hdvpbnRfZLk
JGxQJA3UqH4hGA0d0OrKhdnqZjntrE8CnRQdcj4mPDV1E+YCUs56/7pBDZVnSpOeWU6RXbRMN0cQ
Be8GvLPb8UDYP5dyhK62zsaCezVcCGZWLZxVmcaNSgDi9FeeImOG4WZq9fvmkJhpFCVE+2XJiuhU
jMRSRGluX3ljmzF0cLMjeG8NAhmaVqhESWDqi0/QJNp2urGlJuHwc8ZLA+zf+hfyuUb8VVhTp5F8
JQfkfgCyYL4Eebo2epnEKNxDOnXHsbzidEorrRxvyVdX0fc9oJMKauwWQN9jsSAhcngFHjc1YIA1
EKQ1o3JfLYzRM8tfZiaCPoNCE1oDTQblxDCZ28gCAVsd2y5aLzXbwYk+OOrLQpa8gotjxrmFHxJp
hQz2CPuYz+F0gGm2h34a4I++duBGB2O7VT6PwI3LgJYNNsHcILVGhzX1SlLP5Kg/SIxNpattY/sw
PZhDK+z6mz2AGrRNozfMHzBe2TzbiU3Y3c9gdUFeDdkDELD0eEPSeH//cGsI0WEHLvhzCywp4tso
VlPfBkyIummv9N/SpULohJMUzi/HCcq7j67J68KloGhpZCiOnQ7LbriE6K/wgkcCSoua6qFT/ZZM
a/s3z02Z9fwvoWKIET6DM+QrlNwrfplmIVLxckEYL0XPrUBnm7WGOx9DHXcSzgeBUjR9jV6ogNVq
OXx0IyzUFuvWzC/eN1pxkmDLZ+3Mz+Sr6xRbaFhC6rVAU4z7H9ztblYA04hOlZg/BWxoRQW3ntgw
uGcTCetV+gol2ro08lQFLjInjnCKG077ES/tOhfeb1I/O977+m6g8CaDt9yk+q2GNAGrJoghYyXN
UJzpn5AEwIT/tfq35irfSofe4uTJVWvybZNAU5rM8HRvso9QqRZ2bw7bfArXnZsC5ObmXNka9NdY
XB0ANwHXnVRM2wW7/5996XM9m/t89Iz64dQtQiRjv2+1i+G9T/ZQeRz1kVwITCq+RK1WI9J0Xm+a
Jn5Ck2pPvGIFbOL4mJkCTe5/uVuinxAxV34snySnIHFcd+YiLl3jgZN8l+qKW/uRgDYApBd9cwaN
5QOAlT2gIY86cZl46V5riAOY8L/xBwL5iDqM/K7aagkmNpBWifV4/stgNf66wOjFmbfYyVxP+Z0+
W2keMo9ejgOrjxO3OoxXRsJmRq+1Uas5GJPlGRWzEX/UBdGNZRbeC0YdqVVMkKITeONgcJRvtvtn
dhwzzNEckQ+A0wxb+vZEXNZ1FTEQXWqbtACZ6c6U1mytoaIYp77QH4PEqx5r4KcyFdpc+ZPcpRe7
FPRuuEIyTrtOWz5XveB/X8sgOqW6BngWIYbDrJBRfyYdjNjW+oegm7lswl7nmuEcLS9c2zXwbYPl
49PCdB4hOmRIQIDCFw20QykjEEyxo7xe2QeOZWyEgt59pa5f9KNgryXwnR4ZTkzdJPyYxOkt40Wg
15F9t5XZeMz2aQgzk3BnGeFpGPsadfnRMwgVpST6V46nYT1bBOS0wpVImpiFf/6sWd1Nx6OU+eDI
XKIi1GNC+/xAIF4HaP9FWZDjQK1IXFyTMrwddU5uUbeEm9ZYUJCx0XI2Hq1ahdaW+Sd9T4QRsw7j
NgGj+hVOyh3QZVNODtQLX01vmqAMxzvrqkMVffCS2nmPGwsL3eNN3bzbV/RNInK13VXQR5QnwZ4B
jstVSnO+okafXpFdABng1DyQoLL4kYo4mhZfcNuIPMBab7pn17G1L4AJ+L6AtmAC6db3eAnYixlZ
vRMtqAvNOZhj5bZmGdB94PqffOvqVw4usWe8OKnYUYq5Q1SVrXHrBGxRHTDs/x14eWdjmdaSA8FN
nLnZ9I8g9B4O+CfJLvPV3Cx4s3k+G0wuSinE+/xpOya7mxF6TQ+g/nmyKijXCoOwZGirq112EiaV
UMIMRRkY8WqeVqNMjiruBS+XeOFhela1h+F2/WtC0Un4akeRbN00L6U7oeUTxLC1Ip6KGHSLUFU0
y4hropzRpUC4OYO7byQVE2D2+36oug3pCLUw1jP5k9oDzggr4VvRHsk1/Exb8A33aXQc3oUyk1l7
xh3W9s7XxK4goslPGGrhStaJicXWJgjUhvth8addE3UbY63ZNuTVT6oLUXmi2pjHfaeeqLynIAWN
E9EIy66b1kQywroRZmcAe/9rNlRNwvj354amcleU6PgrFe0YFPrlPL9cRlsrDU51Udp96tH6coYZ
w7b3n7wCYL1AIpWkA7yhKs9BEJzg5Rk02OfpoqKWbF1c+fe+rkqSGs/XVO8zcmXINs19wvqSZvq1
USZVr7394FedRLlmgWrWog7KBHukFQw4fWW26QbdQVv+yEnuq7wQqgFr7p/i+f2CKltHb2IYGV18
E39D7YVMPoaaX07pCUVJO3EoHoTR4k819Jyz74A51J2LinbyAHJCw/TbPa9Z2eP/tT7FKULoCY9j
cV+L2FsswgxpvEFapeXfl/FthcikeRG9HYN8hbU6BRyJwUuxRnp8hz+jRByVaLifBnCh133zlv8W
rw5F2EK1bvZ3PWLT2ASc++Bt0lSlhGF+VT0+38FpncRxToaXI436TVU/fxzzmNm3qqgu4zryANJc
Kowci3BQcroRXOgqLITZSEad/GM1KA3/rLPX87VI7dJ7aJZ+4GQVDho59+msvD1ViLIi3rnMpalA
2kXxk9vqFNBbYWiQ/p70OHuvmnNszhFRfNd0FmqzEotsl8jy/iGWnV9+YnOnOGZjZzmk2jNAPxp5
t70Tnp3Afg+wc5OJEYjQiRTss827nSDHUnkNXZpXXluZtqRVxrbjD1nGOObXPUYq+iIRZObjLPV4
Rx1KG8/p551+Faprt886toRiXYrxbGOBdxSMl3NydAo1OlBjtedADHtP4wKIk8PM/oR26+GVszAm
3vn3QFu6KyCANsUWFQpptQ8+UY5tbQWp+jPQA24aP4bbCgOarLJQBPneBvqQUh2NdbHVpSKVtYFy
BsngQZxFeMGs3NRR0HCBy3dFIFgI8CR7WguEUZ0MQiJzj/kWXzofd1NUJb7IsmTsH1n4tuvf+vY7
Wu65Ot3HZyR23womn7fwUEqSrn1mIS6foutRWZvXDo0Ph/X9C8RRYSb2ZoYUF+jmZbMk6eKYZU5B
ilGLc2VvVQkhAcFqWpdsC3QDjp/HHbr0hUDaiSbfSNaKS9chX+n6+hWe7QoHmA0k8Nt8IWJqLbGZ
242B6yu9M/ymeN9BfQUTav5xNJE6L1PmP9UemTB91PhWwPI9QY75JwCu5W7127G83tv7gq9zCohH
aliqwasKD5TCK+Zpcziv86+F/GhJFRp1Tl4jV9Bugm9ufVf3nE53vadU4zuDh4l3fRofSjyLlDG2
WVJoy5Wch4YjRWfbmUMVmK2yIFMGwNTkytbK9e60FnswWq4W/iwCvxP0sSLuJd7fxG1NVXM+pswh
V+zqLNkeFzHJrveTHnhqlHKPgCodEkAgezHyxhafNTvKrLOAjDX+N1gSmn+QYJ3KvjFJHBMlDj17
zlXAOxWdXbuRWhjvhhvzk4fT6eGFIMurz0u5G3nLhm/WMfimYyda4J7E1NqSn7C0P1o7WttTmfN2
8LcONOzNbLJsU473wVo4mcp8N18lMZrjbIU4AuLvvyLktrcbIQ2IyUQiclWT7B9sthlhekxflQcz
/DGzsHYN1OXyGjm0J0p1R/FkZ0Pq1vTwrKz4aUZtJ4qj+B9t14Zkyv79v8GKb7kYHlnfzkqs74xv
gqfzfLqhl4fYnIcv230WPi2D4BpRH5ir9duh5Q+SXfhTur6bd/lRIKX5KL5mCImCdztcudwSMT4C
prAdyP6ggKGEjVgdZ8uj9QYmGIXDBP2kBpRKvEevLJgFPd/MUd7A5grYYdG2krDfDValUpb46jfS
JNHcCTDVXFbowIYBJCJOE3XStnfzgkzq1fUiNvsrMGt8EJRwql0Fzw9hqWbV8CfdMu8EYxQ6iSwZ
lX1K7STq+Z+grCMqhJp5bQ+M2v+E0wwvl2kxvIFVtveV84BFyZGQ09AWg6Fln5oVsiKAepoFlhJY
d8JNZlvHmslnHplKXoQblJJ7gV7Ap6+3TBAQhxxzqEba8ZykyluVo4kXIbGSMQ7pc4bgz6WBil68
0lgeeKDpaAqzkiwu5jnzcbIPT4urukfPiRff7Hwl2+58L9oKgwIaSQgeqMUP9TciIY+7NEfLLgyS
+8bzeI242ax4tE3vOqhStqqJ1Qwjx1UWsh6Slri2Ai+ZZSzpi/ogaR9xnjj0f1IFFCoWC1TfjkuR
2DLcw1tQaJXgWmRipgY9inAbKWTSnsxvnJ8pK4SGpDcPdV8ppt9eu7TujFuKfESWKv56x8o4aLix
N9nn6a4KcJDUSeLiCteSOQF8aLCKtP8x7P7Hct0ZyEhYQvBWUGmxm3BZQ0SyieaaBe6RJ/oejwVt
UL4b7FEd8zvhHbXsLeAO8jkpQqZoQLHAMIW3NNOQcRlTauPYJ8iZmobZzsPAfoaeY/+bwwRXYheS
u8ndB4EzupuEiUsqrGm4QjxzHwQzr6kujic5IZjIsFt749bXhI0ezmRBEgDuSEioKVaO3QpeSg8/
WPdSTTz7qEhagTyn2rmDnPOnKdQPkdImj4CwrX43pK+WNGdoJ9BnTSguBI5rvPzJTQr7AHrlb5Hx
EuoCcUl2bBpAqDGVy1kTKHY1d9qciiV9qoHLfY9OOIVsOROnIOZR1DjUETSxJONz5l/CgoZ71SEP
325VwQqgu3FUcmu6Obo13fILxjdFKIXPiZZ5Wu5ZEXniFtlJUeKDyLgftxAyzhZEenYKgLZUPR5Y
uxk7/qIWK4kys7u/JJO5IoMmWKblnj/HDoKEsYNpv6T6kpPaC4w/iSVhtbcZP/jHIAMq8X58inPD
vsNVQsuNTflIVZZsYcRyrY8DT6ydgihyx5vpke7OluDkq8Whfy5p9o9/9aDrsDfBxm1r0nIhC3nT
TLuHoUVwHOFHr6A5TvEwkxHce2utuBnyjVvODqNrhFlQiaQxmGu5LVQLY9M7zLhFe222o8DBMfj7
VEKxIM1YFeiXCVWslJpcN1Ayvrpp0aUYsWGLLRBcJqdR95LPRvB3ms7uLMU8V1m/loMTWsyP1zRX
iTFcQQnecmtNA2Xl5OQ/JEHhBpW+YAIIo98RZfyliqnNPjBtraGdpX58UtexAt1fCkMhpsx51jl3
MiRcC8jnjyReMiqGUqqqqjcCjDkiHfciFT1bPt2lEGpHRx8mqjknh7TA5v3ZdHrNTiydGBY/Drbv
PK1LAdGPWdSQFrlgp54MoSOzpZwcTkhuEkbZaLmlznEMQR4gTCIU7qfcSW4Oc5qmOiO1rpGCsqmo
/v2ecLKZNgWJytpSD+TirA59lGaB0+QF2plPEa08u9yFLKS48QyBIShKObXzoF6O6poxso8ksEbA
ug2oUgCgDmbqdgh2Y/56gjaHXufggZSw5KeiA8aWs3xc7s3jrKFi0Y3nlSYjP/h+l6MdGglmX+j8
cgE1mvKv5dPksd8SqdLEexVq17txyzdD2q4HsDtZVwwxu7NhKhQ8lf1nnDxgwx1yxKzChAGzCWV3
CHSsBbNJpux8tvgPP97QFNoVhe1g5KF9tAqiC4qXu/oLoqK5KzCiBZ1ujpKpjR66r5iYC4+AIWj5
BbkvUaOe6uGljQhXiy/QDQyrnEN9kvrpyj9dJzJ6IBKN8b4LOFMXKqCxTde9KI/DViecSa1CxVPY
MQajn1Pt8AnrLOLfb5dIqN+/UyokJUPutp/RC/KlxwL+/T75Lm+OJit08sAZt4ibEKxBZCNP4pLd
ewM8mLMThnjxeTHOXMxtj+Q2RnwcnZ6Dy8PUGNAWe21GycugMH0uDYJ6sm7YwrRDtdxifzsaLqRR
nMWs4eN0kt+qy8groHUPQtrlx+uTRxlzOwsvbx4NikKbDxYfv2njJA77Xoz69ramTfXQr7Ijgt6o
XhCiqUSDL9xAqNbsAFCKtIrvSzvpYf0Gz3W0JkRTDFcfaZNhviQL+aHra7HC/02DHsAoYvF19LcX
0z0gjzi6ph/gzXeihbWmfpzRiq9B3conHKRu196bsX1TkUkau3YrxrwV3we/OiiMpWNzrKwy6VIk
NdIE9KHdVFbSYXi1a5FCpwxlyOCPhm/UOjozp2wkLIM4fJJWX0Q9mfscMn+fW6j2AOoGw/9GAhFP
wKf8Ylz7cbTdErZfimcdtWxeHbkHXENmYyWMsWqSxdmDRceAdYZ/wHNhl/+UhJXpeyGtley/4xVu
UGGRCuTUK8pMebFw3o7z1Fu0y90p2JxBnXl76qA/VNEXZA+4O+eiSDK5ykqLt0zDTmMez9h15K8E
atOFoEpdngORnbXwH3BMlxt8FyxC+gDztiv9Ge7HzDGBxiH6CvG23jbNLDAuoYv+hf5UBK5P2WMm
l2CbBnF7FaS6mgWDpSY4uiMu7EGqJgKsYEaIV8cIjp1kTndhK7hzTuyHxy7zgskYu13d6LngaSYL
/BbMC3T97ZKWvPHrHt8Yy14SvbJt4Ji7mwmxPtSvi0NonR+mrF0oAzwD8PuT+621LjTLkNQBaYZs
j4gr8bFkOPmI9JqemFWd/qC6vKFRFQS9BpXkU2qUlTxQfBOVNbyeVXhb2mNd+4TiUt8uN1bO1/PO
4tIGiumEo5p2/mNqRGDacg3bbr+xl7haFDP3i9nt6ENBN7wPijzhQt7KOIwI/pE5T8tPXwn+Axc0
2bwt5pmZg/H2l/B7FipiJtCzUo0lzy7PvLl4z8zj1nvctv/+opH5TCfFyAc9RJqpX8WU4Y0RmMZN
xbMH3iVk8NZFf368LSh6m91+bxXMZ4uOivh4JE9Rmv/YUmnB3yRd7CucVGhNr0EWOzsbZLto3SnW
h8ke+0jWCo/yJbdp13aKSRI924YiWV7s+1vzImTiSyh0EfnwcqiOZ0jBJJjh29WUFVrMAfPYwews
xM5xccz+7aPQTyU1LB9fwLXmII1umzrfXDGD9xK2PXpdiCNPwlaesEsOwI8cxJ0acZgPHFQhu3MU
LtZiTTxtYvRWd4D3FkxdhzEh2aqOclTRUqx217jDvLFFUWsnoeIdbsTJKyrmeoeQ3F8srI2imbz2
cZyX9VlOl3tJZrQRs0NI8UFt2/e6erPY6LkvKa6PSXjkQI7fBLAaFrp1kjG2h3XZ0touxZNWmsge
u/nokcdPJ9U7+HhPt+lT+rpLJsHUoaZyec9TqlGJbkcfw3p+nn6vfPTWN/rx3VkE9hRZjgywmA2E
AGRTAyL/55mL+j2fhR8nLysJDKTJ0N2pb2cI7xxRg+sh4KOt9IiZ6k1DKlj6bElR0OxqlfqM9lt6
1BJVI5PuDQeHWHfPJ7g9S7mrDxoIGZ/eNNAlw+IDjrDbCPBYQ8EaHB/0nNDMrZOcsO06F9RmgQPa
GWdJE/qELABl8d2XNQB19suFIL3q3XnJL/Ph3sTO/OYPZnrYS3JkbMJNOrZAz3sVbNF1zDe4Q/Do
pNwHqHUGf3Mr6m3Hn0SvNcb1J6eh4mUJXhqIztmxo3NRtmKZ4Z1TcbLlZru76kq7O04X0maoK6dD
FIKFcIrH90FD5BDp/s5I62GTwmljdhi5EwSi6QMqt4bqw3vZ02pNgQ+VBPNPlkZjfj2baiOQtoV3
TH9ySMHTAGGzBIIIn+E6taQlNtw4utV455D0kYNrn5hMIRxMkYpHYCxVaG7LkvotyJyOaNmXB6C6
a4Lnr6FgONlaF4W90RuYOK6A/LCWWyeWbAtyC7AzmsnnVKPVEenjwT/T8L+ys+bG7y00cl5qiVfK
OTg++rcYKcpqYFPkC8bbYuwl77FN+yAVOukdFlDgfFuh0coOQYkNesH/qR8Ge1qePXYmYPQbf/YZ
d4t4IPaAAz/xOGRLDG5/yodYZGmK65JRyWJoNm6J+sS50juW4c4XjNrPqDVeVt1U/E1M1nTO/6j8
DihakqxmtLhWcvkozqbJ2/FS0t47e79NUc5AU1HGktxj7snRS2GSw9u0piMWGEy4kphlkSoYcN3L
HRpmQnT4gO13aGezuMx8g9co6ETtGCRIvXJnBMLp7LDD4DY1I/3QJbvnlGrPGJYtYTkvlUN/7SUW
DlelpAcQkk1T6B56YdQyU2Gr+IdpiczKTHMvA9B5cN8YJPZd5l2r0Fhoc2HSZa8J8RFsj+hf12K9
omaRoPRGtifNvuy/duQh7qL3WTGmAo1urIr+/zdEC2Umiu4Jtm/nd3afYpSN8CAKnDxYdzPjwb4s
G989y8VGLhRBTd85fr63umE2TRyjVPaRLIXHPRCHYvbBC7csidXQfRRc0y+ZcEz1zENIFg2Ug22p
H9nNZCaG9LmmJXr9wbYhZlZtl/Y9TrbjU8GfodpouymbjWq8M/gvlmoA0LpwFyhKGbih9wQ/ELQY
06EGjybR+5mqH2+RSe46mNpEzbOcswD9Y1XbQwimpENJ7B5FNZyMSCsl6cZy9E+4wC0ucmv80Km+
V0jIq5HiD9sggU5YVK45937YsCJv3ss3zXODFrlSp1OdUg2INIHc6Vsi0zkmnc7wf5yiYLXAlAcM
jhdxTC0KBP3uKJYbBpceU9IL981NqnppRgpIDIJndQ4Uq5JcaflIg4BdNMU2hErEhWe7Q+i+ifeb
Xva/kDaJgk6OUj3Hwh5irUC5NyjxOxov65UVwKHK/J3RH87V2y1WtYzqiqlCzaah4FnE0jeyDU19
Y64pOcNc/wInQxzYI1aSr0wQhZ/O+5sTWE4++I5HTW222vxUIvxqpkL/ZJXWMX3jmvCjVGDS8zw9
D9nOX8a+Bual0IyUbOTdT98uGjGVnl+Q3ub9/eFI7hJ2vswddh6RdvP+tLHcplEu3K/8bn1DNFbM
OU5speXUN/3x19gDdtwht0QLXy46IrNnyLr8n2iGLdwpnNHEnJPjcFd9LpBg6+fNa1f8HDAxXcqU
QsupG4y5bNkOwAr6m3bF0/5pOcEBBXTPn1KW1dMq5AdVdGwJSHQGCcTdC1yeduV1AroReu3JcN9s
I4x8dPsM3Y4egVP1St44YTgoz9WwP9Xy/gTLNvkPYBC+taeSjDVY3Uun7J+gmAujZBZbyCnSC/PW
GssT4iu8AkDNWIHcNGn3F/ZrmPxTsJxJieaoByHEdSsyGKoW5PwNPBdr24fBIO7D4nr/JSE2v5DJ
RN4/oCyZnyadQMSwZuwbSLfhXY9tHrVv9637roKMdSeQ6byLjRLopEdzWQjkJw31aygNcMiiAQlg
dgQlO8cy+ikeejgiR8OUq1s11kctVqywkuIgLRppoEghiYHbjR1q39unLgQ3gxrGUVPNw4KKPchc
UhRpQ0WIOPX2hgqPKA5MpSlMVGO7jjY56c67DJpkRa60WSHoedtSTLNe13qnUK7sYxnCFOI2dUv2
Fp8ftfo2bLtoLFezbai2urzHBsUzTP69m/g8iRbQg59+LK0ljS3ZRYrWMq7gGuTVao5leF6fV8Jb
C7HXA5XtjOd37VavjyZpHBtm/9oVOxN7Uz1pzTu2DqhTKIGjGA0Acin1ulD2rR84TG+xIg3IyKoZ
MHHOVIwNl4fpyOyuGm/i6ANmKQh0bq/C4k4xH/d6MI1C6YBy4wGGmiYwWXe5yzbOliBOAU2OM39j
749emjntlAHy471p3TDuVYB7MbQgyFogoh4JgJpn3pnByb9ECagsmQEINdYDQ+lQZTNzec1GoGJJ
MOzMDBAiKHEPo7oIooyPPHhvEJT4jpLifxv9jFjooRnzwkKfCPeWAcD0OWDmdyLNeK1NhwLb1gO9
7rWx/aJPEciXwVGs52prUwqEspyhsG4lyU36sq9S01Hv7WgN7LvBqFevVWODcg4dOc/QNpnvp64T
sxRTv7ZgtN+pJo7E7KGRfHy1PgnLFhQBpHYVOwM8nxsN500yhNxQ1xi+fewxB8veQe+ngG0y9ikj
XXCK+sOkSTDbHJM9jk8R2QQpwi1G5GvSEKmoVYn2GugYoP6UcO+3c1V+Y3ZZlwa9VwJzGftuUKtf
9YpaKmUSP5unqr+VHetsgmyvyI0t4bdDQOnQVbP8/IgMlnBYVRLd+rFmeaP+oaCe6trPHu8h1fkx
SYf2REBnQlKWhQd/YBhJCFMEOSVNsf6L9x6x7xkBul6QzzbISFXRVrXkgtrF/0A9lxWuClrtGfVw
ruZEemwkF6VDvzurLUlODy59vsLGHRfUTG557DAVY8U84vnHEqbz0wvXab4wReDjDh0kIG2nT5+1
Kd4Kjsxgz/G0KVFofc5Qfe3jevZBJc1LVJrUSUh504m3oCR2NgLN3iNMCq/eZhX80lra2xbpnLTD
cxiccZBWWtfP+Q8ToPAEwvRjkvDcsyY4oUHsv9VvM1YMtDyF2foTn2UXEVDsylIciqnIyA+nFnYh
LFW8OxGbft7n5jQxiAwNu0/O6rgjPPn/YC4+vrd/SsRXxWwLr2IQTN80m9uBZ5W6hOYPP0Z7mFZL
e/Kebn8umZYWQpLmFTE/gOweQaVWgSNMG1YkXU+y40b7QN+Flut1YAbsg4Ww7GjQ3ofEnKH/S9C1
3jZCGbTgi+zMssqkWWxZi5Xpd9itrHobctUoBjcxw2uRIrMF5NjE3012e11YD27BZ1c1LJSYKdrD
VY1E3ZTtPQs7/61cgMt6icbn/7VYNSa/VZ3cy1eKn5WBwK/58XZFG3soqvJsEXgaZAI6PEJgCEsM
oqFBbE+7AuA9QNL0wk5p3clRSrMzTTC73xQpRjpk0MJrZ0/VBAF2dxOD3mGadygG7peX+HYoT6nL
ju+eeaFlPQfA7qMT65w4EUm2AiAd6lkp+eNdjA1xoPqWrR995tKCEkfn7yvcI73kpuH1sNMaGBPq
qf52EEVQeWerNiwWCmMzu3Mw0o8JxrjnqP2QntA3nl2tt3N3aJPMwLdP0NhJEjORMYwAlOH0ZKZe
6jeX10XUSSBzjGgn8Kbzyn1s4Wxw5UmZfjJve0W7p6HOjjZO0kKgUkEhywSNVFQkyiw52k8hVPnz
ZeHQ+LxywoJ7lKQpggFRBs1znsrroo+uOxw/m4gLQz0FX9c5LZ54dutD75dm9eTyMKPQ6ESe2pmS
lMFB2og8HsWqA3pj2g23vmB/WVp/MNg2Zj6nUm78SOpR3j5aTC2kxMvMJojc0k4ufwrqHnxmLV4x
arPpKCcp8ASUO9nasp/KlrS4VBVkJkKZvty0DR8+QwXg+sbYqXbxBJiA6M39CfI3QRQXCYWUEFz/
/91qsbkk6OQoCuPt7ZOYCkxSBCvZWqSQEPBgU0T3QsOXOIC735CQM7x+22sDGZxlYtcH1b/Frlq4
oGWQOtEvvM0YWh57eu4+B/3oQV9krl/JQ/MjTQ3iD3iIzdCWZFsBkq5Wa2VwdhFXVmPFiCnNpZhS
VaqUqTc/nonf0F/zj5X55LlEPrQA/YRdNzEWhONKOftziMyk8BXEaGQwNLR68fkEk7fyUq5XLYD2
t386bA/Br1BoK83lS3F8cEvww8VwmtxxgwLR0h0kgrPSpONS7s3TkDEhPlm9xEMdWilUxP0uDogB
4yD0J7cGwixNMDyMbKCJp3CVUZzcoHjzaFXajhLIuAxqObQhr4je0hr0cv8u0LtNDjVStTZ2Q/Je
Umo44cnkvyWybiBNEr7doiClRdF5SYxOam7H0O7jjMjnJRPcIz7Q03Ih701PRd7bXsSRyvHdMRFd
WVjPGoskhuMSRcmLDByohGYKlWb+UW76SeNRcyT0NMWz3192r0Z7Xoe11HZB0xzfguEquDH1Zpk6
S0VdlJMisGWFx6eepTUUKWpNADA9Es9n1s/DsPY4jwCtIi7APEcZwaO9195O/W+2HhMnkSYQXrz8
fAYxhpe3wtbfMx8bzy4FF+v01K0IfqtiAIxe3BD1Ac03/jE9Dd1q0IJ85o4g1/u/CN4DK/l/yvKO
aaoDAM474mK0uNVL7gdz7d7kYiBLOCPP5W58OF+l4GbHn1v1ban9d3J55xVk9UwNYUVUuiuMZCaK
ROft6Nqzsz/92Qgwov2X5hSjKTPjWrD8nUklLls3FKDfZl7g/BuaARdQ3eK0XD2eymJjQmDiAxmh
aqKCbTj56ePlq5/BiKfMvEjwwZjBXZuk/C2ukquR887Lqbhh2E/c4TL9eXcnKEzOWYKSr3Ajcsgw
SHLFA/CD/Xibk7+8I/V99tTAToycgquMAR30w0w+Ivth/1HTd9ENutpf4sH/tw27FIq0j0p5vG+b
RJVV5tuC6sHcYCsJXiEzTNlKbAYbIMeyxZVjObFj9LwVI5YCl/sHow3VNxr8kpLVY6LlcJRLAYgd
sd0Gl1zOqG8aqXYDEkG8j0JHTmI5oLmIQIy7sEgcMKEoS2A6BJe37BT7aSSlBHkCN8Q9xQF76uoo
L+ZW8/2B95Cpl4ReMr8Ap0Kw4ZVWkunmbCxVCUiP4mGNhRdKUZU2AjEDHZpSM8CnrqF+TyhtUOkC
QfvrFkMC37aUKN98ZzeQXHuOU/ZtI+M9UN7i3bfWPQe3nsds7JAUT9ATABtafe3nmQ8Oc57AugvJ
JYk3VXuZomdlMK65rXLd0hwhyRMumDp0la56a+AWIl77bMHgsPR8mXTtjgu5qWSV8hwLmpZdEta4
L4Dk2YiRXTXpAnzp6wI59nsG6HqCdrHr7sEevGABH0sFSfWIsWx+s1yDywhMtEpJDmRsD0Qib0I7
ii69lhU0XGcbxYEPQBnC0HUvFdP7eHoUopmm3TfLP8Jgsxl7EXgDxhAoLgaFObRGi5cKObJuxY0A
xHG3RVjZNtdjXHupnTE5YMP+eaEIfhffGZLLKpLSw9Y1jrJNWDACslec6vI3ERVYYxCq6zvHytWg
ztBYF4B1KF+r1K89z3R80hQqhnqYqAvFw5a3Ca6gORlZToWT3QfCKCYJM6jyTlRCdn9gD84FP5QS
Wjvp8rfR+Fm48EufUB8sk+xw0Hrgc5p9sjwrYa9ha+lq5qW9Yh96WLr/C8IqJXV/KJCZfWjEedVA
47KXWxisyKWDiELNzUSkt2/ldIryEKPYmyEn1OqEc8jiZ24gfvUy02EOQz0GEUeWRPUYtz2cWklr
M/BC/UzYmtkM6fV1OncnOnls+UQK506LT8ysmOqp8Qc1sM+VnxVpEu8nmXMkkr/cXV41r7SGrx7b
EEYVBrnDJCyv1N9lKLu2yWNsZnjTGNSc/NKyzxNAHTqmWravGKTaw8Kx1GI9QaAtjEF4Z/sx1+/j
5DOwAz0hh1Pl536I5m6ngfUEWEvzfDf/CxawtVhFv8/gZEL5/B+neNcNEnuZJpdjtMZrcea5Hy2e
PAA0JdtF+hznGKhMrsWaNFSUaoh/L7toHf4RAdHQa1YQBJxIQtgfkS16mVE0gtMCd24W/I8patTt
R+N0L0tJGilw2IBqrbVaYnCuiC/EXEJ/Oc/AyIDf+3+Ag8GUcPme1OyB6erKdxya4OnVhB2y2MId
ja+nMzUV8CXIRMAAKApknjLaF09uTxqNUXNrgkD/DCwbBqKAo+LY61+4V8Pmny8KOVtxNpTgZN1U
8OlZS0/FqVziZUdhx9IgWde/5E28rI5SMaYglFZj7IgdPnmVnc3o7FudYNNa3t0dCbzVurKxb6+o
x75SCWWq092+XYMOrS0Nr+AaGxvcf0wiJ7oE7JySGaEtZ2A+5+ESSGc3gP6BS5JmNWwNAl6wuRFS
M9vCzCGiRf64EvLz4oTRnUUNlf0x5E2qiwr6z9q2ZIRYD4ohueLdz7MSjtcOa1clSLY2VkH70Tnd
ZMpYtSZrniKq9U7reQ18Qi4dHek5NS4HfUOqzov4MsUCVMNriSXTUXvtfwed5y2/+lfg13nXwJRR
MbKUf2QtDBbvk2suB1rRESMA8xbSnc++ZuYQu93be6tbysx72ZMqF+FfeUlmqYwWjidN4PNHLY5G
uLsfUGxeF4tlfSLTQolppNBonkR7jUfi10HHKXtQ8QjANMoJp2+vtpvPz6CYP0cRIKtaSsEOcLxj
l5QQRUcim5BpYdPXppqbTt1mmKHy3ivzqaXZ5Mpj8TbacldJX8/cmwqH4tt9nBgciTv7g893kpAg
yN7v7eOuuKkYk1HgAUmAgX/koJYh9TzfLyimbYyDgSTKwhpYnVEAmc4Se1RwPADvQsbKIBkCpf+x
eSfb9b4c/psd3RsL/YEbTWhKN/kXQlF+JTgqTaThgnu/Nu1rT2ao/0hnWCByifRzqAMgFZVrq40u
WMYHw+8kf9zEvFiUdwgoTGFt5OXVmzuU5zm2e4u2HrI6utlxqiLFkpnMwFXYlNxGo8Lh/LzzXGgv
3+8VCO9Q69gbTQ8I04g2gleVasaKAnfRTtr5hFf4JfiGmzfJnRJujGdk52Nyimu3dFQasJXroZJr
XTITfSlCbxjS3q6j51HOleA5srb7RreAMtiDjvhu+SH6ryZ24SM8dvb1kSerwEGVu55TqGNXQBzl
oVfoo6dga8Ks1Yq3zyQWWhW4xV9zErSpWaTlRQOob6ykDZHy4MJQo+lhhbXTZPV3p025qRQ6iCBP
etfqkqc0Y88LbvjY69PFUr8zhglKmMJeCnrZlLnWTM41+LMrSsZ93ZIGlO2tEHS43IXDyAuj6k1R
PhQly/cZTvhfnXkjO6KFekkQSHOrETQn2a39aCbpxgjObtSYedQoK1zlhFLppieQsd9tD74w+mo6
nGcY09Tz8fvT+9J9CVk4A46mmd+IRUKVDYCknRjZ0mpWphFDutu6YuJMZXq6NyL2yhJsYFTUgF5d
XCqgqv1F+4Dh5i0WLo51oIEHiP2U5fVA52RJ6UNw83bGwcMCaOPjNpGzklStoeajtdGPhdRS8BaZ
DjcmTmWgoX79hhY+mWrFjCpAVqvZZJm+5R59ndBQauwW60cyh8lg41i+XIJun9vWi3/bcO9k1MnH
HiFx/iE0nJCNAFPLPRnfgZvWX7O4u4blvCOsziUaJFygr8KkEE3iNcvaYtGyXUW3lj3hbo57bM5q
0qhd1biBBw8BwlD8BZm6a3EjPM+LGI6B4ISKDsnhsy+u07SX/AWlF3Pw5ZwaudaXi74X4HZWMew5
nqhNXUznvJQfyEeaytUAEGlDvpilxxq2VSXL70fRZ6wZtgzSrEVK/7qItkldktYb1EHUO1gzJ7pf
eV4FWeDIRSZHMvsH7QGA3oTG2ON09dobYoWE3CgtBNhK3Od/An7jLGM2q+Q9/KOsXJglqXfWCkhm
xxQ5O0oD12J11MIPQsuxjMIGUyaaK78YHnQ3zhyikEZ390QkOUXBxqxrPC2fg35+aTPUqV9RTixc
M1elwP11meuJ+6VXIzrRGX+nnUAtmV8YpyHC3QIdk+xNCFo+a+ESSs21or5BmLLVRcxQi0G3K21G
oNfHAMrzLVtVfNm5OtlYBSngcMwmjSm+glX5Mh8ZOgw5sGZ1ieW9c2oX/Lmq2N+uZgdWkQOKeaUs
7beQ3KDfhsVS0Mv3hTq0r16x1RsAYExtIrcJE63b40ijcesgq5GQdN8+/LaLGh7ne9KIpnyS0ij3
5bF4qCHwE0qZPfFfpml4Xy3hPWphX/SQQkxi/2jUz2G7ufOWEEcYWcwfW0N6BGdoro4ajIxbvClD
MK2M3K3UymSMXRoyCRcDKbJELnt6NW36QULlpfLczF1jWsNnomIm4H1CmnzMdI0BDxH2THKHTHTB
WKrgniBDPdrANnJ67w8/BnijXd0oCnlFu0cg+tknOp6ndBxcoa+xQvBFhIrK26iGkUfDJuGrOaoJ
HxeE81wXB4ZLdoDPJvJfmjx1WGScT0LYxGytkYOL7GD9bGrALbJpZfM3DemvkORNWkXmJVMuaoXV
2NWZN6WI95Q8gIQwQC+AD9AC0x9S1fsKN8Svt4duTZee/6W5hj6kds/p6yWAJqLjAmoVi4sE1tDJ
Av+UCUlc251Qd7r7+mEvcQVLJuoQF0OtehjIoghTsmK9CBvqyuYGER3WdMIiKoMPfcn9krIATjhI
myOoWVTs5VHxvs+vsPCu37fuh+ZEVOV264p4VUVj/se/fCN5l+CNQUmLRUVp7GWStsZUWn0qyDhk
KyK5cWgalFElesRx/aymszACqKJCb7mgPQPlS/KbLJXjfDuOkJhJIDYPv1gYSyytHfLKRN8IZJsm
3+3tbMs4ZmBeZT1SyHvseG6JzGUJz1XIK98JSk/WLjQ/Qyju/MGxlrKwovYi7/Hy9EqM0CvVTyeK
ofxS50aBh4H8DtIv7R2fhIgnvwSzxz0Lxbm1WScJvQdsETgZjmQ6BQ21vfm0iJuXRUjpZF7FiixK
doqsaKtIMJIIPJraSK+aAai6kA8ghYJaGy7sYfKfgp0J12h5oHoidBNiiktNWRAtSdWviO9Xocwv
7F7Y/pUVBYVJSfzC8Texkg2ziuRpkUdqtzJZmB17f0hmEYKdMTWKq2hfn72UI1L68hsAPnofJBhQ
QuEq7JBaschEn8UNkMlvCA4qmSl+Fr70cNYH263Y5v4oUf6MZdrO9Hu4c6rAOwCXNfXXnvW/A4N2
Bpncu/W4ztTCGYJCTF4sSq7Xx4psvJlpunN4iBGXjHA25lV2WDdT3HTqdNo778N3DxFVLfbkx69f
W9sHyku/VXb/CdDAF8CVz7RtCzzUo9r4odvBKhIj31FMA8uJlKUvK8pgKwjFSAhjs5BZIBHX3DJO
JfPlZxmgBDzg2GHlS2z4J+kS13y2n6/rpnJXtbt5gnhsk2cPUjaipLz8dUBPbxNIKnsydV8qinsg
qNchIk6xBIaF+1yEnlRCTi5VuSJgkkVMUYDInqb7W+vg2fiCmtnP0j384ZeZ12mYhE3QkgxFY2Pl
Dm7a2L1aNNQdg9NTHJlFYYHcLJxuvCcWPco4ehzNhyXMok0wSy1YflI8QMskIP2TGNbK1+m0seAD
wBJM6PaPzdKLflOfyUBmhGcKzZUmC2TsltxIWUsW6ENULXkimqpenPm0C2bP5qNzbAxvd7tmzf3m
AzRKIA+65BmisA3cgbd4NACD2LgmXlGFcgihUAehelel7AOggfZT0hjoqPZ14BTpfe0hf/hUiNl1
8jzoCCgQysSGf3D0YBaEHjIxqtEouHvizcbZOUMqnk5HtxhNxFph8Bo5jz8sLkKEA0tgQ4/oXNh6
Gy+34E3OD0hINybquq+tL7XFgVYGF/aWSsUIhyj8p5rKPUzk7LfqF38l4zOp0c4VQTBu2pmssA+i
bGl8i4YHirYGpFpW1BPwAksnt84mv18pAXFa9nA9DVhzUXTg7ZHbk95f5QaWhJJ/f9WmVb8bglL2
AT2XlrVrl+EXfuy2DlQHxKcv3gGp1ZlkUG1Rbu9D1C/BG1G3UEIGyYYEnF8iXDk7vAwPqhkEkT+D
f26SngMozsph6bevgrrEjGeDry4X3LzF9Viox3cG8Kgb+qLySNOOqAI9g73zmnbTovKvujej8moy
1YrDLlGiQxgpzX1P28CLISorNSKFwZn5P79iwwhKWmBvUad0lV0uYJ0jT0iv0a8DYqaG+oBX84wc
e4h40Cv3dMjKgA2kSEiZ/2Jdet3Jp1gOAApuantDNxUBHrJd+9vqnGetrFMBeaxsp8iJNhtx8/cH
s9SJH7TruHAL3nPjpndCN7G3vGfGhs7QtSohmfwFifHJgxwnSmvEkMjaEgWPBGp+qpRS9+dyPDiV
PS3mHEE37m2GaySpI7YHNQY00s3IW2eMPu7Vep4CkC84pGTO0rjc3kf5Y3aFDtaq6DAdI2AXrIha
O7Bs4KlwxbRG2g5gZZOy8XtGYu0Tb/74s0OOpqew0nJHzNJpmYArZkkuKVeu9AxS+VKNugAl/K6a
PSGWvpkxGBJAGa6QlSoXmjBzJFHy6G9PVxj1fXPcVOj4T3cZkCoYcjaNtDKUu9cgMe7UpuKWq4xL
JnDPQlybknWQJX0HiEZlevRT0HGV4XeY5dinVJLr5z+T0Q+ZqcgUDOkbd5/pTtDKiYBdm5qD4iUc
ZTEV6fLXfLyNyYLqIH12cIj2Dm34wkwdo9b5Y7saR6ortatSQ0hH7Z0nU5/AqQA6GWgxYRnq1e5h
rVwqrvC6Ffs5GDkCJq9FRoGWbzEMb2+zUHvZFnIVLjTXtrmTlCretRMWyABADAfhJD4MdxvZ4NVZ
lWwdRiI2i7jzJ+osY+M1h6x10OSYxPZy3HMRFDewpdPBRtJPFuTVFPJwt0OcYy+Pck1yh/Ize0lv
m+TsNDw/LYvmPS9dZ9va2q+4MW9e5K6QIEaBaVDG/bFLighP8hhk70G1qQbJpzhSGkZizwMCqv8Z
Z92ENjmuS6XSKoyEwZK81EDyKEn87utdLkrMnwybuzHudH6stopEc1StA2j5NdZDYqWPiTgZb5rR
dHPeGUVcT/ealJKm8VAObMT/kavX53YiTnMZxZr21KId9MpUuJM3dEFSIu1idzjO6LU81BPERhQ3
r6/e61zh/pwfNbgQlW33z/CwrsSbBVSEQo2JQ65iDIyicWDUvD2elIMzlWXzqXgobCYFlbcwvhGN
jT1zm69dU9Ltw+xEzP+XOlo4nV3wVDt3eI9l5d6GY7U+IzGPV08icXTHqhAA46nlJWjt7FNx12O2
wxUHamvNMTql0yj0XHm/3EHUNZN6HUerQwfeOZcM5MP24KSVpBl3lfH1rppSqe/OVKwbvnAdWNwy
m1brj4i/Jz+6RGxoq6ta0TlrnRg0bHjTfDTVb+nevUY4crkmsC55M3sfd4xOvrJytSNBp/cg/lT8
9lIh5Gri/TTLEcVMc3QQP/wxDlXaLt2rXfkiPHLHsRgmJD4AdReSGQg18ZfsTQtr+ORRrODnrGc/
zHuyDVM3xHsd5JoccSRKOksq2xIXxHs+6qOCKdGdc838/UNgEczM4NBvfMOJau1BVPK9X05md2oe
dspo4iNF81X6SPO4gaV8L00elQUnH/kZ0bmA72stCwQKIEWr+nFigFkEmVk4Y2ok7mxFVgiFQeKH
joPUEPYLXHN01OF5Pn4h5CfmscwBXG85Sp1UvwcDX25rW4rkazMvKGosa9580iZ/4aEHd0+nZO5t
YlQ6iNM7QvTTbFBN3n5GOpxVO6RgZ6nMZQcNolQgcgd5AmYqrW+B4m+Hwgq3VdgeDue7EIEVNlZI
BGHKeZlvZfyUGLSR0K6ULqXSxAGJd7NhuPZx9X3h3//l9XA+2AYaL9uOkzOCGPu4JRyRUMznl2sE
8usnkTGSDl67olIKZqTXKwFvpeGv1LcMUyTFst/m/VU5hXlAwaKhe8liHf09uqIJMs7mLkPiV56c
rb6yhlFfHZ2kspQFAkfrDhshGgTRPgTJ3ZVd7ltSgfWNoKAJUfrnAXArHOkbsNMEN31L9OmgXKiw
JUoEWYhhu/IXH+wOMFGeqrcutYsNPlNRqWTkdQHGNoXFBb3DZb+Mt3WafjGeltLr4JudIqP2dpEs
t3HnhXv2txWPDuC+bG1mvduPeZe6FG00PziEhF/qYVSjt3pwkHCptMFOZmCDo3WeWEUGTwHxu9yN
BkZHJ4cBJ1s824+hDZunp3HSvf3kX1urwqDhPUfjLCMLF+3BTSfCW/YjA/9K6WTQocNbr/F6oIdN
BdFHF3z/ylQJ3ClY41s8aGmZlxnNMyHLde2uYpBpb0hmeMw8dbrSSGhjSjcroxxhK4KK46T1vbpd
eW53R6scEULZBG975PgGSeCctcsT5ycTno0biHuZcEubLIHr4Nvzb/j4E2Yegmi4Er+Rp1Lo2gb2
H6aWVtkRC0kT2JVDBWjVWeXI0aP9yCBue/njrJFGXx/57+87mHqPp1v9l5N8i+4Wi4hClfR7UMR8
jM0v+w6+4iHv3d/+KMcf0mN3nHsJfU2JMBwkVp8YrYFK9GVIsEyrsCimZ4oqc/IVxFY3mde+8Blt
8Ctq5D9eIqWsrvvhmPnVPcChVrdD8h4ga1NLXbZtA5z1b8V+57/sS+ZOfECpBkSg44GiXIoVdMNR
qlNZ10uX7uIqAbTlY1scGBS0Wk/3w7R86SaGMhwuyggfR6cM/u+kEl3HeOaUT6nPKaPOrjujTeZu
LeWyvPJGhXlNkeWB1ldR2GCrBXyDiZ0hw8b1fOl2kUPjY7Vmtk8J7Ws458G/w5wxJEljC4HCVwGJ
RAf9z1KMz9gQUj8lvhMfZh6rBOV3a1vjHUuSCIgPmkVGVyLQrS90BBaycgbBdW1T5icn19vtbPgG
aVDK5izLc92h4sGyz2HEnzxS5YGjAhp6p0hIxSFyMpZ3XpXsgDAk44oAK2XyBHvcomDOcsGCKHP4
11P0iDTepnlFLbeVl5rzjUEfZ+C7tz5MAQ952NKdcAbj3fgUsNs428F3LNVF9C1zdIzdaSR8vdei
QzDRCvUxK0VTRBYkD2afuAl1kfy3hgAV8/CKkHNFdGgPHpK0KJIeS+AvOJxCXDu/dR7q1oVXCXVY
IjnjOP0p2p6Ud2a7znN5+bux5FfYnldV5zhcmT3EW7aSgDaLucTgl+Wqd/NOMLLgpAqbFHs2QMfX
PXqLzsfl/J7c7/UyCSb4Km+cofCuusvGPdDh1iXtwnb8B0Bs7YH0FNAbQlPXAfIqYdH5t+cxlupa
8YmvvKna1Aewk2hsgal53oFWCGFP32EPp1z3x07luyY13dl5fKhxVGy+bFOhPv9G8wDUykDxCWMB
JxX7k4yaVfwsBlmynLpwLoVxI+bUH3B82fB+PHAf2CvyxJn06c0Js2dAr9YE5fBULpVN+y7u8IOY
gsPzX62wn72kc7xQtMjQCoe8IvrEDcUjOH+761mh5ziTWf8gnl8gt9553uou38qizaxF6ebG3jsT
d68ertphKjAr4xqNHlXqQcHxD5vhiCPiFDwjucVG14Wkt9581xestbOESk3zKldzrNsgSaFXeEAb
ZVHkdWFu3p7X3xrUdoL28YQLvCPCdrYVtpDcB2i/Hc6NhaEF/s1vcXpcugALu5em3NzecMfctflS
kpeK9ivLklQZMqKlPnFPcvH2FJvmadbd4OHWZLnpfI0LbCtw6G4fxm/V4/iEyyvatcgxAAMnzt4E
tKVvjxeVzj7RgwZZ8vKD0rCiKE8SZiYPghmYnNM5TzfEwJRIVRS99WwnYdV78jpIMjOOh8GqiawQ
eLikgyWxD3gPh9fqdUCVLrJw5YGiW1hHPyygN/myIzas2tFPq/+apIKpxdL5vaA1SpNYZlAJojHN
SHC818j74Re+ceJB7bOuYIpGCbwHFedxHp4SOd2kx/M6lCkT8kMVO/1kMMaQKd43/cv5P3GvQp9Y
79/OLvExlWULdW16sPPPtZSCc19xmMF2PwMzOoicNoL0cLl28mGqv8MXylrabr33UKJ4PS90oUsg
NUYmcecRZUdGaMFQ53fwWTao+q/xbQ7AGgKRjXlKwoNSUPgsmmq9Lw70RjZoGT98Gekg8Sre+2GT
jRyZRyrnAyMWzGNDOliqqXA277YpHQQ6hIRZUGIzGrfn8AMOL0k1aLsURBy1sWQzOz8ese8TKj1z
UyXKUzR+TspXIoYgjh5qSU0S0rfjCqA66ZadEupTPWaToe6hBwQlHs3V7di7Yvs5oLUcXoDVjBOo
s56gNy6kq5PmGWeAPcbfuYLk7RuSr+w5YRfbKGGaO56tC0aDyW7e916J2aEQD90UIQlq7JeExFDy
yzG9hnfiwV/Tawiqp6EA5kX88+yjGWd8kz82T8WYA1LPHyGFFWEdqI/yEaBRXixrWlOSLBAy/xtw
tOdB5nM05GbQBWTgSEBhNDIoYSJbUVqCgVojHrmowuBZo8XbuT6FxdVHAQ78P+dlVrtFLw2JnJFB
ZPna3T+ikUosNzWe8OUoF0rtmF5BFSbnhu7wWXr5lB0Zp8536jm0KaTUnTPt00qKAPJeMo6V8WQ6
vOBrG3We2zCWsz1ZRFThb353z03w3FCcGrpUV0wsn7O9mCk4mO11W6OYdGKOBIKpI/wqMKiGwP0Z
kfkceyKbEeTpVyMd4QRqpdFAQXO4EvShmKQiOSVNSZHkjXUyCT4lNXxHCnywrEVJ/Smi4YIe+dpx
5NHz4dc7DXXnD3miSwcKc2p43GARVfAOaEq4ZuQ/RCfecH0ou1Fbeoc+ligjn5+p4eCIjilJrh7Z
FfwUyrXVny2sy8PfaKrOCCEJKOgAZI8efiaVJi3uZpqlC75tKpgkreHz6vrjxkMHbGXoCQzVQ4jf
yYJybhK5cywxzzXkLS0AEX3XbMm+pIbdkfo0nuwZr88TRJO4SVENovAkgF/VOgWnd3aGJu2gVD8m
Rg2R/iJkmJyjiW8QVlOKuuvZ1gWZ5C66/BqzGy7a4gz5ukRfJKjT9ZgN00TGvn3K0HWWOTCJQrTp
FdmGcwz+eCEhdT6gTXqVHsSCk/0VHeVCFbMQSk9M4uS2s57KeNuHWF87mo4TcPbdlD67OyCsnHtj
3N12q4KWq9aa9aAe0ZuVgUFw5CQHC1OuuIRVd3N+v7nLkj48Cfv7fLQQnSEwYTailXiTGJdLecvV
jLNKtG5ujusooohv+CrnB8FCtW1QrDD9Av/YmIUptVUM5T6DIQBUg6IUgxc6k2PTeaKqSxuA1/G3
HLbbikJZbCTI4gS1VQGiJs0cIRZFr13X8F9R/wuY2VBtJLuT9Nxz4OZQkBJYcsA6ytwFWVJEPyce
LDrZV79pl0+gDcBY4SqxkLQPcsvlXlZkJICsryzGcrgBc0i6w6/4+H0uNZsH/pjiGxoSxlh729Jv
bOjGZRt+sTq+jH1v1dev9hsMiXuXddFTwIFBX1bgq79HofhoD0DrMQc/jCa7zp17aLJUT67wh50W
+JAOkSrDlylpxs3lgv36aJ4MvsvcSJFZZeDwGpl1fE6kd/Ibg5tvATFKyVEpibNEqmI+dWV4vxc3
KTapbmO8ryWcaihBsFxV3sEb5lzm6N3qKyO2UahNqzGbSgjo46AEWWZllkhb23xqns68OhbO/Cch
EEtHQ1cjBV+5/ymoogHp9zSNrVtXL/4xWUOQXLLyXb0h0lJHPSbVpi75unjGfJWTZOw2NUudgHky
P9o7e20UDa/oLTV2mxf8sadXat47cmzk/O12dxwEqpPuvHPAzOqB/nbcC8NMoTRZHfY738q5ODB2
Crm9+SwIqDxvVFOzAdX0JY8MkuxE5OGWanESXN+YGBgnFx0YVl/+hNQ5wjkThwMhIiKIx84UmlaB
5fo7tCYjUJtq+hQg3bSRpwbSn9MGp+8FiDe1fG+ep3CsgSd+t8xnHs+z5wfrOTkp3vGrz/rDhxOk
UzTdw+UbCcCR1ndwkAcYnzLfIpNhoRLlQ/+tM6EHL7Ub9B4e4z1lWHVqbXfi+bpsIgJd+IxLEP7l
/5Eu/Rh0A0MewGVuZ4wYSttfeTE57VfsWDJAx1u7VDgsY4LiOxnX+5cip4TsGu3ObT0s2KCRw7Gy
MbUnc0/HmRj9jMiVaiF3m89HczyeJS+PWE3kaVQKpiKEKyBtTjdr1L65ryp9JB6UIMNU9M/wwfj0
jtJpvsMpJRFE+57W3vEqY5srwqb/yiRULEFp3WAm9ak+aoSbElu85duGW26treJA7cMf0PAWyiRm
DFBQJtevmodi74HXZFuekdIPLKWP0MGTJbD1Niu/92DM8NBYmaCiIkb+FbxjTFqfFajhdMN/Z89E
I6T4DGRyIAepibNmMJFhJ3kIoCXJPGmUFsjra798lSojV7xMXAAhTJesH6zPkvwwIMgCx98ByISR
xn6mqGAMT/v+TKmuc9OKj302y8D1s8HAj7jic9Yw7zCN6wqY92yhHVkle7QhGSY3TI5uXFEzE7r9
X+t7x0gcsM+TT9A8+6OYKk02j4CwXYBG3fPzlLnPUKQHJ+DMJRzbJoH5m2b1ZzC+/uISfOB7hguh
KjqmZelgswNShyRxKtGOEBwtyTurIWrSiPBxw98G6eFGPkg1ECpezix/bgauvB3lx7252BdAtCqS
svg9DQW+8bxXocg9I8A=
`pragma protect end_protected
