��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2i�>�|���B��,<��\ ��W�~��O�?��K�މ�ͳ�^�}9l�}�X���*��Q'����Q�R[������ ���������iʔ�4+F�',9�88����q���h��Vv:4�<���90Rϳč���	ȭ�U7���&,!��K�8
.cև5��%����WD�zF�*Hjx��ؔU_�?�	S/��]�w�$\S~�S���<������}�r����h�>�~wHi�)"�UM��U�w~m���1� ��^qx��&	9����b}� �{�Q�oĽ!�7%�ָ�I��9�}j��Y�z�x���o�Iŋ��6+F�N d��o�L���X�=�S�]q����EòM-�{����B߇��T�O�r�h�۫��/9x �����p��'Q	��W��-�P=�ɬ	Gb#7>]o��%0��Ɋ�^|J�L�-n-����@��;���g6��˜i+�r�`׊��e=�ud��&X��s寁x���#�j4� �x-�ڪ��9��	���ɀ��`��K�K���q]���|X'Q�I� O
S#�L�S������ŗ��hd$�tQVw+X5}ab�YQ��p}N�>8~�u��&�.��Gl-�M<>��\�p��ŷ���	�Xs�06�p�YcW�a"�:�,W񠉡[Y��c����<��m��kreT#T�EłS ���'a�oP�y'c�
P4�����\�����"x9�o��脛@~�9�+0���JS�T�b�ê%e]^GG3˫C��+80�J�aV[nw�C�R�W�2��r�Wl�EiW���)��[����Q�'Dc�j��x�+��}c����-����j�����l����a4T2����a:��=9b*�Ίp�hEOb�T�!�dЁ@�|�NU��vs�qpiH� Ux�(|׵����=�s��ۢSf��]�m�~4쑟� ��B�'{MȾE������X7g���M����
�VD��K:i����F�0�:�l.���QmH��SP�Dڮz�? �!�.����,xq���/y�ȥ�6���a��2�r�I���Y'Sb�c������z�6D��?4�wxO����� p_���F�T�ފ���u0Z;�)�
bm�oѿI�=�ʂ�K�)%��Q$l�d��=�r���M8Kw����)�����vB�Ѳ&���}`�j�� s�_�Gw(��'Ir����/yB[ç���6l�����QZ��|��E���bur*?f{%��l��7?�D��k�F6Ͷ�ּ�8>1q��B�7����_]�w����V����|��y6y��0= lH磨ϕ��̞hɴ�7���r��������+������?�u��o�7��}�ǻ(�A����u�L �BƧsR�ݾɩ�z�u�KjF:]˔hy�-Ϝ� ���M��	O]l�")6���1�;�O|E?lݠ��}`{@� JLktٛn4�W���#�J�8�~g�e�$J���i����w��&�y���e�H�5_!���E���*������	���[ɨi;�:��~ϝI����\]rDd2��7s� 3~;�H�<�ڗ�"&y0�G��{^!�тw��'��F0��+���_�+a��=ᒆW��v;����Z9�dsJ�������
�ъV�`B�F����7,�;�L�"���4�i���I~&'m)�����
>J~�Q��.�W���!������jA��J��qD1��<G[W�����x��o؞�����N��f<Ҧ���z�	�a13���w�I��zZ�����m��G|�6E����Q3j�:�$�e�6w�*~ЀM�-�2�\����]��6��#�獯 "�79G���߬㩩�r�-�jAU����[L#�k��UH|��_�h��.�<���䎹����L���p�1ݲ�k4ӥ�^b�(1���態�A"g��G��D�pzR:(��6�;�p�8On�U�*k�\�`��C�����r�h4
�-(�h�	�mE��_��ݝTfZ��ʚ߬�L�LA ���hH�z����<|�)�-�6�.�9�F���n��zU��<�(B5�o0,#���q��E�^8��\T��-��~��8��޺��.� jN�*��[���a�/ĲJ#أ�Ԭ�eZ�M��7R����m���"�`��	^��ʖ�u�q���|F>��USd�s��c;
�C�H��Ք*�,zޢ�1畴�E.�Hk�s�]lݾ�v���B�	����ˋ�V�v�b��	����@��K���WQ炼��GI>����qێD�ܾ�I�eC{�ұ|\��8�K���Dh�]�R	�J��@�>�������W��y�Đ���G��Z�Io�Y_�r������&%�U�W�e����m?��2�wG��m���r�J��󰼣��(u�� NJ�\�Jp���oֵ�����y��|�zO;��*<�z�14�I�s�"@@��5D�E�b��ᰦ]��w�y��iN�(���Y0��M`Gj����Qo�8���5����ꖭ���b8S�ߺ/���68<;���e��,���m+PBD�́A�1��!��Ѿ�׭<���y���7Y�Ig��8�wɑ���t��`��S���I�x��b��~7�~-P���ξ\Ȱ����������h���usC�!!%���ֆ�9y�:yH	��7
��Kg3�N)x��/�g�~��0�0�yj ��v�?W�_��?���c��H�o��6J�@��1�<{&y��Aj��>?�̯1YG�
�U+3h���Q�l�u�&�__K�&A��tܶ�L�s����lb���0xF@�-f �Η��L�
�k��e@�UM3m�N7��&��]�P���5DwC�*�S;Nȝ�Ug�9�߮GҌ�{�yˁ��W
��w������b�/���hQ�LC\)�)?ZSB����#��t�k�<iv�!����
2����YȾw���{�
�+��*J)��!Ǣ4/4w�>h@6F��gBi�VVi�"�ɑ]n�7c�D����&�fx�F�9�H9��b>~V��C`zˑ�p��Yzoy�̄�R6��OM!��U�g�p�a9��Fpr`Q��]�_)J߷M:.a�uc��|�]��q&Nt(���IP_�]y'�Ä?��
EED���wy6&�g5'`O~�||�ۋ�3��>�S(Z��&_��JU
�dfؠ�WE�8ib*_t��Z�D�1X�]��MFrl�e���x�����g�X�BCu1���U�L�葭�݇ZfP����H
��؂��X�3��*�,>h �D_��c�ý��,�B{�E�����2��}L�P�2ܤM�ع�~�J��{\L�����7��	�:\�qڇ��,��Kp�g����eń��I�M���Q�j���e`Ew�CM��kIf��*�j�>�P���L�3�#��<EPB����ֹ] �Qo��/�l��\��X ��VpD�k��5���^�[ű���8�zb�
��ycV��q\L����5�ׄ;��]Y�ޙܼ1�O��,�]V���]�����/��5��K��3���}N#Du~S&D3a?6�!�?Յ��:7N >�0�[�{g��,_�yb��7������^|�5��]:�Rى�u+�ݷ��nT��P)<�1��-���p5͍ L��.���g��������s"��[W* *L#Cч�$@ڨ ��ܼJ���YII�Vo�3�E�H�$��uC̏����[f�.H�\��k��
�v��-�"bq�����p�3ӗ�{�������=��.U7�\8?-��}<�3$>��@�.�����G��C�S�|Kn�{^j2���;6YHG�uǔ&�$�0?z��j�%lu:���?�\xr:I��IW�Q��?���/u��c��V�����>��?ŋjg�}���mn�	�l~g�a�?c�V�BX��H�<TKLqhuD?ӴH��=��
7A�:g����ź��ǒ(��&F/�B<d:��'��)�tv6��n��5�=r�o�����
/��1���`�Ƌ�.�B��+��!�����5�E-`bZ&�8��&h�����7z��i����*=Ntت���&7�6ʁ�2-�~vn�/]�}}w�p��@ܗ��n�L�~����Ts=_�_;�v�}�V M}�{q���"D�����ʚ����7�+��(w�Ut�/Ӻ�C�#c�A���]X��/z��v���_���'<u�<!��U�oC�BNNrfA�J�+���j�M���Gޤ�Cy�*C�_��V�^�:�Y������W��0[��U���EEY��j^D^]�3�E�Ij"�k�ie�s�+�V�%V6C�˩��,�^�����#�X��1I��թ��į˾
%_��<��
D�m9/d=�#�YE�h	����[�W��n�͹1�
uroT�}���J0:⩖Ԕb�D��D^߽�0{��y/?Â5������=�b~~u숸��>_(���� ,����5�n�q�uv�X�����p�$qP~Z�9VN����U����d����?&\1B?C�~u]Ӓ��^��PZ�v�֤�~NzNvC�w�l��Nws�L?�"8^��-����Kw3�p`i�����> QB�x��ۡ~��Ia��5d�P�*�i��!�h}d`�����R��A���A��d�5��u�	��| ���vnm�&�>�Qa��z�:1g��N�+WIjl�����B�>��[��R0V�p�jJYϳMW��-dt�8t�-�~�'�+�f�.}��_���^�8��Ě@crN|=����g}`����T/N�$�|�(�X���\Y*�!����Q^��P�o�X�����A��=00���-�ٽ��`����ц!){~5B���{M��q��حI_�+�����*��M�+ww^�ր�n�]������$㶤лhCD��L�Oh��⚱�*��-,���)�|���y�^<L���~U���[��oƥ4�aF���H�)FO�p��>'8{��xW�ݗ!#>�7�י���Uq���E^�Y�l���$.��L�ќ�Ê���@�>e���e�v�&��c0[ش����:�̲�_����	�f�Ӕ	އ�nӘŗ�s�_��g���K.�ڟ��W[��f_U�g���f!��]��: (\�|ҖӍ%$�QI~��
����8���d��.��t g���� "����/����V�偖Aé�<����Xk� ��8!l�pȹ����=���o[̖E	�?�F��U,�'��XJK�\�]�cbؽ7Y�K�9��g�v�������D\CΒ���n1k&SqO��������#y�/l	!��'�C�-�w�"�O��;� "�F�]{i�JCq�~�O��_E���Ӄ��Z�e��GLU,R��8@7�9 �^�m���>6��kO���?e狍Ѝ�w�T`Ӡm�0����oH`m=\	hs�Y9���߻�.�i�ch�*b�@���l���.�JLv, l��;ל;����!8�4tu�������ݳI"qzj���ܜ�J�T� �&���`����rn��Ϗ˄<0��G��0��m�<E����'���ni��^�溏É#�Hg�
��4ѳC��r@,`����"V�/��X\���htm�0���4_ǡ>2{u	ˢ��(RBP-� Ml�F-�r���i�7��H"��u�����)�Γ+��0�)��mOP������F�'t	��;��F\����pu)BX���&�OJ�c�� �����{?����`��L+V�6|��u.�]:P*��9�r�z��_��vtS#���5lD��LDZ��A#�������~�϶����e�tכ�4M T_�H0�>Q�S���͔:r�U�(�,��j��Σ��?��7^���b�����3����R>�z$1[���N9��T���Wgg���ͽ��=�ʑ²mi��俛�&#��Q���R���DR��>�<�/�"D�b7��}�]Z8t�:I;���v-c\�HT��$A`�y NsGs6��_����[�l�nc��UC�V&�-"�;mF9�w�t��\+��3�s�?3y�j��DQ�`�A��q�ʂ-rU�����Wb���Ș2�EF�x@Q��R�B�B���	}�-W����@��cdL��gH��)Lm!�P@ÚD�����:��]��F��������L�d8Xފ�+���q�	`8
��޶�����T,���Bd\��%����m������uL�N,Q�혌�W�l��:M�>x(�Q/M��G5t�kNޜU�i���A�cd�����P�$p_I�������O/�c�s��c�k�t$$�m��8�*o�T�G�rZ�Y��D�R�낧�~=����C�[:ꕔ���mVP[Q�3���N����&ѽ�!V�g��@S�w��|/l����Ha���V��1�^�}��5��bvF_��}~�*�A�.��qe�pЯWL<o��gJ&j|~K��	�?_[ӳ�(D�oL���K�����@X/�ٕt�K_8/�U�i�%��Ȓ��5�j*�:��@�"-�b�Vj�����M�"G�΍`S2��F-o�
(��c��9N0O��>#���Z~i�O�.���#e��_E�$��+�*��/�-�5�K!�;�"�-�'�[g��E�X�y�3���G�-�!B}s���>���m��NF&�[-��]qC(X��+���q�Ȕ��Fb<��SDӆV��M�a�9PE<��mO*w{���EO�>��\h�lk� ��h�L�K��1��ނ�ߓg{$�/��a>�i�#+�5���(�ױZC�)�$�ןY���S�o��-m��g���G�+:�D��!FDEVqA����6�k��c]5�cY=+��f�>���D�8��DŔx���{%V��j�`O$7�_Qj6��M\����D,%f=5��[˵��^;�Qŗ
����"�tdZ��V�1+�ޣ_��ćj%��v�W@z�����[�,&���J��g�d����(�l���=���>F��TD*�����&����fuӜ/4aۚtq٤�",�8�y����!d�
Ӌ�ҹ��qї�A?�A��X�4mp_t9��T��@�Z�̨�ތ�r_��i��F@b���E��Q֚C2����-���3Gy�VOkT(�/sg{T4w�<�@�����yD~:~è��h�{���&W��v4�IW6ޕI�~� ���wE�>Q�A�o-	����d�m�J�N����q��:5L^�m`wAj�7�������g�=���HH���;W�['cQ���WE�]�@�:�5N��5�V��W.�?i��{��[Z�Є���������	&��P�wƩ=%;MPC���|f�κ�"�rw��� �ܦ��9���ty���QW�J3�u�Մq.�{&29�<�( ,���ܰq�&
D��Iy�F���l�Z�L.zw\�I5���UI\t��R� nw�\�$��l�De쮥��8V4?����b�ݪ���>%�D.[�	��Q��F1�Բ� V/h#�"�A'd\0�
�;jv%��iJ\�5�S�|�&������y���ek��F����<U�<�ݦVzưͺj��8\�@s#��е��xV��fK^ڨk�xVj���tQ�^�D����#���Vur�Aީ��V1���L\E�7�|�pw(�a��5�4#c�I��Z���)�1��b��'CW�D��Q�<&�E)�CO�����ӒA3V�rt@1�
]���a|�� /�r���|<��CU�b�~U���Jx�
j� :���lX��v�h}�
�W�0���nE\8�w�h/�Yw��q͈��+&/.��v��U�P����*Ţ!d����Ӳv���@�ŘL�34M��G�V��fa@���PS�u�He
g�V[!f���Ju.�����ѕ�T�[�F��<�V�\S�A�]�[��:ĭ�D=��釧o��eӗ�3�ڶx�6��M��\gD��64 ��{�H��x�ӝ� �Y%9^R\�`M%���K7��#T5�W��]7����&�h�F0�L�]���Z����u} p=y7y;8TtF�&x�
�M���'X=
�Mn0GsfϬ���q�<� ]#H�^��8D��(R:)ܑ�ze7�x�GH���i���e+��I`�53�,f9��TY���!�p��<A�5б~�I�։��b�gsϤ���@z+��X��jۘ9��F��PY��!�Ζ��8"hk�ǭ�򸠴���^���x���S4�㯢]�ۼ"�R�Q������Q�u�;���2ĭEB�"oXxi�_JVQv$i|�P�Т�6U�c��_߻���gr�5B	�c�VЈ�VD��6������&�cJ
,)]xI:�%�y�>�V8�I-�X}C+�㟅4eA�#e��.�ԭ��" ��A;����M��✼*��Q����h�\<Ę	�]�l����g�������V��@���ژ}-�F+�d='�����,�r*� �6\�4�k/����x2�V���9ti�伋��,`� �Z%7$�V���nһ�����^.�;�+*�Ӳ��������'L�x�Gb��Ѵ���OV2~P�oWw!8'S�`�ܾYA�ߣ+������X�<&�DК��?�m��ց�~4a(��]J��V�@�f���9��k��׫�b��j#�
_FG6JQ������6��d�q��ws�Eo6X������$��#q;7L���@��/��/L��u4�o��
cnn�_�3�o��[��Y��"#�W�0�CZsL��á`6sK�/�����`M��v�･X���e�H��x���L�ǅ��o[��JL�Ȩ��`��!);�N&.��e8x8�f��)�Q(��/^�lk�,=�c�g'�pr�Z���j�sI ���q[º���Mם?$���=%�6b�^�"Zq̏�w"$��Jz)��瞃$����#�'2���u.��L�Kӡׁ�b�o���?��	!���D��K*V�~l_ȝ��N�涹8���� ��'��#A�6A�»IG�K�~D�L�=#�ĊE�Nh���.W����k�1�G%�F~�8+C+YG�w<��a�.x� m�X�����K@NI|���B�f�w��M�����ڤ� U�p9��{Q}ZE���!��վ?�G�6b�߸G*#͑�����L
������A>��E1�6�k�0���j��DU�@�j]8��Υj}�#��s�ݙK6���{_M� 8�kk���)*��/]p�z� ^���
)aH^u!o� �Y���!͋/@���ܯ��.�suX� k��*/�&�u0�2P,'��=��Y�>�<�iH���n[}|c�[�nE�Kq�5i�9�a�4��&M�	6ٰ6����(�7аe��l;F�7�9���W&���-�ƶ\ ���Y���5:�p�p��$�ډ6��%�3(���ڪCi��N�r#R�-��ڲr$��s���ǀ]����J\�_�R0g��:N� ;�kت/h$�wq����nA�����%�L�
����!�& ٟy|������P�3�㋱V��3��d`���;ú�O�t�7`S�v9�_��z�]���P�7h:sT[U�m���Y�V�u�}Y�aP��uj�fe�lγ'�{���)�ֈ��8��Zв8��O	�J�ы�..�i��kO?�N�Q>����H�-
�� ��2k�~s��A��h�=��t�GG��0B[�e��ߗ3/�G���4�;�:ѿgy�YV��۷��X��;�Z�D�X4!J2�J�hB~��ǐ�>JH���=u���/�)��q3Ā���$7�4�\/F��"��΂�9��q�`�U2�l(A�l�������`��RG�a,��VӠ��D!��o0���T� ���xn֤<郪�d#a��t�	S����D�Sa7Qռ�R,���G�"�� ����Q��V.=GYx��� �V��P�a�6�{��D`ז�]�x�aW��&�R[)����0�_������h6�Owk���*�1&c�s�k�#ms�H�l�!�\"�thx��O��M;�b�?�QFgI���u�*�؏j����i��{'h���iu�v�eS.
��KĽ���@��m1����Ֆ�1c)�0�\
�k�t�����gR{����p��j���觖�ݮ� ��5B�e��x�ru����m�c�#Ϻ[ȶ��G�A�o��='�(5U�c*��h�"���7)#����ZQ4#��B�r	Zo��} h`';_�}��gc��wr%��o���{>IN����%�>�D�G�û�,%w'Q~FԊ�愬������2���A��v����ˌ� �N�5��0��s��1���Z�\2Q�;#@���2�;�9FF��5��mO��ܖu�ڠ��ӎT���A,@��~�z$q
� �-�2G��B��sl�ቩg1�S	h��.
*��(�6pؽ���9M0���a�� ><�F��LR�'^�pd�� �Ѣk\Y��Qj���f?I0�R��ޣ�6���e���H\yp��A�9e������(����ͪ�Տ"��&Ȣ�W�`؀��C�b��#fd�%I{����3-�������6jW���� �܀\�97J�棥���+�'������d_�D��B�ʯl��&,����۫���s ����"	���zT�Q?lv�;0}&�=kP�ߤ3r�"�+�)����g�כ����}�y�r�WN�Q�G��D�,�P��2����l�2��o��G)�2
hoH������r��y��9�n�nR%�����$�so�Z��VfY��� ^g��A�G� �,�j���u�A�c��+M޸QLD�Ø�W�t���J����&�-۶����L�vk�V�y�t�SfV�����j�q[��A�
P�z����M�dƙk�B'��jW;t	,7l�E�t�n�����|�b��FxS�Ub�����b���x�Q-(�ږ�d�F��. �/r!_<4�t�͠��s'g3�㌔w9��Ac�!<ݢ�Y��{>�nj}"�vL���,Y�=�2�2ݼ��v�D��!����Nr@��ح;���c��G���:���T��˻+ƾ�P�`�����B��}�x5=��V������N8�����j�<y݁�XJe95T�w����	UF��x؈� �������lT0Z����5��|�LZ�"�5淥e	{����X�,�4�|d�*aB❬��N����o-��D��\y����(x&T7��I~T�@ͯ�!� ��4k��?@�L�%�ڰwѼ�콣.M��t�����~�����Է;�&�ӳ��d�%i��c�E0C��[�Qs�h��Re[���0䳀�SM��\
�����Y���}6ׯ�:�K�]lN#j�z[��l����G��6I�1� ���d�Q�NjK>���4D���e�6����+�h����p�7h*��#p8T����j �q��F��D0�qS9�z��y(\|X��Gq��G��G��0/�3.<�Jr@�l����WǦsE(>�kVjlq���\��s��s�L��w����U�B��&�F���(2JS���n��gzMS��u��/\ �ط��)�����~��CsLk�QD�8�~5��vD��w(gB-,􍃏UF81'o'�����$ŏ�TJ��������˨�xS~�o�홶:���S��r��&^t��?��*�>�"���t&��Mp�m"Q��3��r����ma7N���o���B����������^�%]kq����ehO���/_���B�j}�E&��^!�f�p�f�NJ}y��2��]'Ggc	mWMQ����yѿa��tة�gX�Y$�����ҹ/ ���4&��tX@�����H������;[�<e&0NX�i~��?ϧᐷO�<w[����^��nP��3�vÏ"9?w|9(���=�[l.�rOO��UW�h�*��{4����z�dDmCƓT���xO��*[O��թ%'@i�,r��\����%�Mp�wB�����=.d�ã� Q0�l���]v=�R����:���<@���f^��EE����cJJ}y� Px"9�A��F�gTNů#H/�FWٻE�h$k��,@��V�/��7Hs/s�O��)�O���\u��� W��7MB}���B|'���%��mm�̓�W@�%*��-�E����� �M��E�.fD&��2���߁�!hRy:6��M�G�I�^#h�o�*�/(����	^��Q#v��P�Iu���=JaU{tzC�;�\_ z"���Y����Ҕ�F\�N�`��.��S�,��^��~�_(&���@N������''��~�Ӥkߘ)���>�bǜ�+�-rP ���=���qB��P-��_���j�W�o�Q�(�pF86DBc�j��35F��r\�$��]sJ��%2���ۛm���N(�"�����`�3��kI�wS����Lg6�#����q�a�j*�%͜4��;V�@���\Jj�q�Z�q���%�� ��]մ#4cȎ��J��:b��ؗa���W��q��(�Z����4��[�&���+�3� %�B̪����FG���uǯ�'�	�`Eͱ�K�8w�H?gf������m`��ؑ�׳=ǚ�S�K���\��"�䎖�����u9=����P��%�+�=� m��:U����/�
u�����̜��w	;ς�:����G?`���LnإR}=]����҃��RO��4�%��[5J�q���&��V��#2�8u�ܺM��LG��Gt'ڠ�\�O)l"�3�l��+)j���zp�H+o �{(�Ϲ}Qi"���B�x�-ً�{�wx&J�I�SX��W/�y�[����{�.��k6Z{�J���n��*�si
����@��C@~��(�7�*���Ό:�����7ϗ���t�]X�A��?�b��y9�S��l��S��.)�`�3��+'\�Wb�WngC��O��	�sb�6�H��F���A0���.<��5����Q~yq]��o	��3������EW�|���}�ۋ
v�N��Ca��2��X������tn�D�!:ԊCm�9#`}�B�Ӵ�����u�7�R)��ħ����3���:-"n.����q6���9�!���k|H�}'�:ڜ*pd�R=����-8\��y��h+ ��Qm�Ŀ$�Nt �x�"�'1���|��4�ǜ�G*��JtY��aU��Ƣ]*0�؞SK���A<��u����&mMy���˨��N�i/�s$�$��]�����_��,Q��pgJ��>?����������n��p�apIvP/��&�J�>����N��ug��\YRv#�_�}����
,^]���4
����o�X����-�Ps�ô���IR���3�]*8c���Q��î*���l�Ҹ���$�)pYL���K񄱋4Ǧ;��UQ��pC֦�����3��%��g5a�ik(n���<sEe��/5Rke�ҸB�eZ��^���m��&�6�m6��d[z�2gR�=reS0(3X�y��Q�� 4Ҭ]Ց����<��ܺ��Yj#�[>/���h����X�cf� u���.#䖊����T{��Η�
�M�;��]EZ�e^�C18M��D��}�(�������0�n%�v̌�M{T���]k!��!�����M&ߙ���_�a߁����>��0��N.pAD.�5W����| ZO�q��x$_y<ҟ+�V
of�w`$�]o�"]*���'O��tK"ħ�
���J�h�	Ig�� �Y�m�C�댄:|�
�؋Jp���i 	(�T�=����J2��4�߆����s��c�q^��!�M88�t���v��T�Eqq������h��A��u�J��8'r[�ܳ!C�T5,�}ݒia]�I,�"kӞ��hp�m����";An
�����ո��L�m#��1��:����q�9,�R��qOsC�0��;�z~$�c�yG��B}?؊O&��83�@>��ٮ���Iw�7v��}Z�z���>���L��*�د�|��]����}���Y(v}/�
R����5*�!��7��v�����@���!i�r��E�I4�(�ؕ�}�M ��9�$�~_��V�	/��*�c��"��ϊ���)OԱ)��uQ7]9�L��ڎa�ԩ�xp����ǋ�#Vݴ╛զ���;�Iy��1��?�t���m�c���GOE�)��e ��^ac�W��ǥ��b���\%�K��o�i�L?B\�6]S�rV��ɾv{C�����޷��oB,��д_�i�fơ!��5�	�ǚ"ʎ*�#|!�Ǽ=���]�")��{|Vd�ƭ�1#��� �N'5�8��T%��uxb#�����h*��6X��}{R|e�?�4�Y�
*�g��0s�FV�8�ĪA��ɩ�*�ϤFI7�&R����+w`!|W�V�؛!۰��Wy�E��ܕ��e��c�g�f�v�N�ٍF�.�M����qYo"�L��1q4⿴���-x
�I@��of��i�8U��0��0�r� i��[��=�i�)|p��s�}��O}m9Tĭ�Z�G����"=���}Z�YR�r`=�BP�2��dw������x�kM��(�t?�m�'*_ϑ�O���:��v��uT�G���C��7����@�Q����fi�ۺ��B÷̢���y7]�w�wc�+��������"k�n��s;^�2�|w"�渽IP^x��u7j�"������8�"x3&��l�6����K�>��%h���*�R�b��B�}�,��{��i�g�趱������'��H���ɒ0|O>#r�B&��������#���b߶2&�c��
4��:i����~��&������?q�8`��%�Zl��>��e�$%�?�V��T)�.��@E�l����d�َDt��dni�T��)�TWӊ��}ڡ�F���~��G�ݿ�7	���mm��~ϖH9��=��5^谲Lbc5�<e�a3V�5�1=pE���'2i�7�B�rm�VP5�8�;�A|��+��v4o���3�H���g>�D"�|��j�A%��Ru����#�z4�����v-;o��y<@�G�ά^��r�I��Y�����gQ����%��}׬>#�=����hxƙôG�IC}k�{�ym�Sr�� ������=�)�U���>:���[g�yǁ"��Y#U[k�E� ���e#��^K/Yr�����:լ�P�q��KS<�]*_�!�P�튿ȁ]���zɄ�P�O��|�-Z.Z��!i��%�&�V��!�=3�2H>�}x <�x�k���2b���JOl���~���t[���P�������`K��6�|¼6�s�BV�[���,O�"C9Q[vưa�!gp���9~j��g�Ǹ��/��'�4��F�2x�N~C��1x��u��Nc|�m��۵�;K�at��� q�X����X57�.��n�I���S�Y� �D�*��+L�WP�(~*��V(�q�.Ե�൙Z_��[on�cv��6��ϱʊ7<��g�I_����Y��]ED�{��_�N���KNv���.)/��ou;�D�p{�'6X���p17�H��Ƀ,Y&��n< ���U�Rա��/��h�`��p�V��ר�N�4q�Ňx41e.^o
��)̾w��,Þ�v0U��\�Og�'�Խ�����m��:�FW��	S���%���]nYkw����#��_�sM\8#�Q�5vD1}�������N�.ž�*	��Zݑ	0�X�-҆�@�p tJ4��dۄv=+�C@ű�?��W�Y�t	>�̤#�4#�Ʊ�M4�ߞDx���("ɯS$f$����Jf��o
1R�6_"k��,7	W��w/��o6��6�yWRv �c�*���f�K� ���G1Mb�!ﬕ�˓:������h1R�z�B��Qg�#�Y ��<���ϕ��M��"����.����s�-#�IkW�.�.�~�T�C���
�C#�#_E��<!��;Fy(�^rl Ek��T�$:�e����ą�R�rjs��
�_C��kX#P�>f4�3{Mk���Y��C�"���\O�e�I�'���bvsm
ߊ8�d+Y$��J�uヤ+6���H�;������l���H���V��=�ч{҃(���-�`T<%f������G����A(x�B�:1w��1xx���Tn���x��V��979)ړܣ=4�l�܃� ���k�,���^��IżdX��n�����MB}�֊�IF#(iאo�ț�RuEj�>Dz��45�����5�n=���tR���a�#��:��� ��c8 "��V��;�����CXip�h�_I�������[�㾒/b�}E���_�}�maċ�6l�0u�}k1���FpV�B'��9�J�j�����;)�_����4	C��"��Ϝ�	����ɱ\+S����!�ȅ7�*���=ٍŰ�ύ��Eo��73c4�uA��)ʺ��(�ۋ!�W����<!�?������d���j�t_^����NB��isYL�ڇz��u��3����pS��B�v�L��K�"�v=ETXT%@a~*r���_g�������U�k�I�����!X`�b\���hZ�/?'��F�m}�-���s� >CU��7�x]������XY�M���&�.ne�zI����dtS�}M�wr���F_dS�c�1ܳ�w۾����"�Ԓ��r+b�����h�-�r�������X��g�
��|6#�8����[Zh��?��b��h'u�������1�����
��U��-�*�7�{JPzt�/E���ͫQ)Ψd������5~U��E %E`A���H�ݭ,/�p�I2�z���z���Hj����y�'�P`m2V����د� ��G���d�A�P��t�z{^�|Ǫ3�n�x0�,�y�k�=6¾h�CW\7��\�x�@�X
��:�#.i"��^��!8 ,J,�!�5)���+R:(x�;ג���^^Y���%v~��g�)fW����R�:��}G��#U�"��S������t���d��,W�]glP<���fh�g���O�W��,�̦��Q�+{kγlu�5\�=	 c�o|:r�&�Ǉ]��k��J���e���mg��tXWq�iw�-nb��	����*s=ʷ�� y�fH��t��!}�'��':�@/���\��o�/�0	��d���feS�P_wPd�ڡS�=����GB!Bb���.�P�����)���@>�Qqs.U��5�\�Ԉ�ꆭǘ�p�����CǆI��������|WQ	���/���
 B�����Ob;� �'@YM���Z�����,n�^�èz=u*il�������Ȁ*Ґ��x$���찾r,p��o}YA�έ-����(-���~��8��j�	�������!j(�|�!����Q���ᡬ4ǬC��8i���$n��?q��z`�GE��{͊l�7�Q9�n�Ƴ����@S�&�g(���������|7p�����/Th�3�Z"۫��4&��JD���QG��� �9&=\.�(�
��c�SP/G;����0)��[�u�S~P+N�;��:V�-���d5 ����+H��,/%�EN9��Q�ʕ9obf��&���ݻ��<C��G�A��$�^�[������\�I-�ߢ�&[2�¤0;,��9�=���<O9闑��Vo����߂gE%��� �w�7�w�"1����O�,�+�P�yN��k7m��Ņ=O^�9l	�>�4�K�R�ԋ�	�苨�ͭ���k��{�(+���;�ԓǛ99�Тt��[������BMۈ���T�sV+�&p�8_>}�+�����nr�Z;ɉ�亢@y�؆M8�.g�w�/wa�[=kh��8I�>1/�^���0A��?.�g6�S1�v���@�c�]�tc� [d�7v.gu��KW]fg�����{F��m';��id#9ɖ>r��q���#x��zl������"97��du�)�{�J����n��#*F2�[F8�/K�d���8��ְu����h�bMC���P_:nN/nzH�c(g���=AC���	ִ>���7����O�w��f�nn�~��Q$�Sna�db��-a�O��Ro����󭱚���j��a��%&?}-��Y��0�QE�I3,�kԄMC%��,�2����0 �3o\��z�Q�\#?�I'?�	�����K���ܡqӆ����%~)#���֔2�~���M.������t#�b���)y�x�f����f���$Cm԰ �䃬[Z��&c]�vdA[�K��r�)~�s?y�ғ���*s�
5z���MN�{9u���Y�t�A�r�?O��Q9}�_����)��E2b�\",�:k� <@�I�/�&G�eV#�Wo�f1��QJ�i�U������u��Ϊ_�M8N����R/�������<m����o���5���� "�BG���'@�K�#��Ͱ,���꠸��6��ow����8�ІJ����a)bO\FV�ߢ�~Z��=���9Z�k,<���U�ݚ�wV�S(���k
��N4{�z�2װ�w�`��DJ{Y��ltͨ�>�xjɘߊV�L���OD�6"!Bi�T���B#�þ�#N���To���R���	&{�4dQ�X\^�4�xW��-�U*p0Q��M^��I��2����\��Gَ�].�}:�eW�E?�����Rma��*�ϧ���^m��+���=�gQ�,����x���*\��<��+fw+1
�uf�b�Z�t)�5g�wsX�������L��pP���kG��o�ɪ�nC����؆;����>@���.���網ޖ�J��/P�5hM�cɠ:��������`zO}���J������A�P��E����RL���뭾+�
9�8דH��
��5ĺoJ��g�����KC�V�*J�Н3t m��1��_��O'�����s3�fѬ��M�/OO��ʟa��G�!h�����R��5�Wޓ�,L�bḷ��� �L�=/�-�Ss�,��Ҷ�F ��Q�8����D)8��20rKb�CP����I��>_$"���e�KD<�kNl��,�����Y�I�Z�O[_�;o9�`\=�dg�����%" ���X:[7%�]Z@����^�{�j�E�a�{庙�)v0�E��R�r6��|����({�b,�|�G0n(�����%	��Z~�N��Ok5�:x{`xP	YT$��(�G�)K�w�MOe.�OGRC���{�8g!5�[����S>Ӕ\ǽ*�ι5��J^`8Eq!�B�++!��@���i���}Jé_h�wc=�z��9ɰ*B
�I����}_I�zg�`+���.�ᎌ!짅s�q�K�,�ªD��hG9�L�:� ����H3ݦ�L����/9i�V}M_n ��|Z��kl��V8��4�5��<�I��O���r#.4۾U.ӳ|�����ߘ��_�\�X����t8�J�g�_�F^��-iB��H��ŋ��B
���L���Z�}�9w��U�w��z�q>�e.ߑ�C̿g�D8��8�$\^o�e��l���d������6��0A�ޅŐt@��LmY�����i��ג^:�R�J5+��RE]d|�^���Ԡ��y
�e�0�M���陫�����8�1�^��q7L��9��I�r����HV2�1щ6��1��Q�y�ښ�lQW��w�N~�<������m%���������ʪ���#sڔ}`�/~�7�^9��[i7�2f�{҂�j��&hΑ$J���-`[�ѺNB4����_���S�^Ē��p����AJ����5���}| �̣/�H�Z!�w�9��UO�Jb�.�����*��r��>�1���_"�[�}�BA���M��A�ao�?c� �&n(.�\����b���Gv��8F������m(NB}�ʹ5���f���p�E�P�m@�(���6�w�h|Liެ�f��4��|����+�H�n�X,��y���1'M{H�k�?X�S�eu�ݩ�$D��%�G����ތ�Tq67f�8��|�{Q��N��{u��JPa�?ൗFf�����1�����H���~�d��[�Dx�ء�o�O�M�u��>����|W���鱁����d��Ĩ��ӜԴi�{o��&�)�Xh�Y��(8��(ȌN�0|��p	%Wɳ�*�G7I���4NSWJ��!�ɼ��2�b�
x��1�,,kl��D����>:_�q��0�	����VN_R��@$�5�K��kz�긹+���������C-ω-��%#͓o�׈I�dO�jD���Uq��������.]B���"��$MǼ��3�Ⱦ����+���Wz4a F��'B�������Y��νhk�I^�u6���W�#E�m���bia�}�2}%u��e�d�� w�:��殝a�2ub�J_:%0��a ��<�Kd�{6�*������ z��$�A����.@{	�6,Q��Pz�^-	t`G�z���\�5�2ҩ��y!��l�ĕl[�A�̝"�	�D�0�b��#�bI3�cg�q����2#R.\�C���w���|%ŚT�>�d�Ι�M~�c��n9Ȩ���r���}��"C�/���ܼ~�#��o-�KJe ����$#�fl��
�C	�Z��{�����w��	Gz��\eq���3�#[X�:7p�����M�r�\n���'�l����7����f��H<b#�Mc[���eʔ/�&^8=��V�6eS��(���F��pOwT7�b�&�����n=�����)����;zo&�K�1��JW�|��i�}�?k/�� *�v|Q�Q�����Fh�=VU�e��Y4a��+Z�m"�%�M[�	�Ơ� ���y�z�I����zG�*K�w�ȣ�E໣M������crb;��g��z���c��j���H��o?=���N2�;k�B��w��O=@E	�a	��������Q�743���
��/��̸��5����?ʧ��C�/�VF�M�G+��*����va(r��^\�x��ݱ?�Xj�t�drE�h�c��%�v&�Nx��z*0�m�'��4��������U�����E-I$�5��]��P�4��~�V� ��F�cP��c�;��0���@��țƂ~�@�e�w5�bhyh���+q>󠝱3v|���v3���p<Y����M���5v�R`�0L�h���bJ(�p�������БƁj1Y���,��Ņ�.���V�;�=�Ť��(H���G({�@RO�����kBf��e�NW��PM�l�8�8(�$�T؇WLbF���V��@�cJ�1=b��(���j��ݑ 5�?�"G�=JT�d���lb_��&i�<V�@>s��d ��K��|~h��`��kyķ;�_��zy�=��]u��a ��K�Srb�������R�o!�$p��Pk��q�+���o$ YݰA|=�����c&�Z�>h���P,��u&�0T�M#������TN�^m���\j	���S3�ς���*417V�j����-�����kS-(88ZSC��ՍA�#9��[�W�2SJ�6������}@l��Ho�i6��Ā��#� $RTVO?�J�l�b��I�.8�a�ȿ��2����۰��-��;�U豰-Q�[b!�X?E�G�^A	+��@/��˞M���q �d�FvƦ<T�1��Y� q�����N.�c��T@���x��J���<In^����� ��)�x��W:�Ʋhl��Iw�u���"c
�u��Am��3/��OɝX���)ۏ�:��Ҭہ�E��<�z��2�^�B��+_��� �T<���ܐ���9gsP:�W�6Yߏit|��Ѡrͭ��)�/2��&d�y-�3���C���q��S��9��q�S�u�Zk�7�t�{�S4��6���' ��)#�)*M1�����}Iڭr=7}��sw�Sj 8����9�6�nrA�r���s#�x��V��c�������C)k�T,>Μ��E��7R҄?�Ney���!0�]�*�G����2Ǐ��%P��1�2�N�����^�A���u�6�c�	���4I0>�~� 9�����P#���w�}�[�@�zɴ�h-n3��y���^>C�{bn�@���s!PC5!;�"��i�&t�Q������ι.��t?�r�;+���ݧ $ϙ0C'���^69��s����I�K�}K�dm��E�H�3����mk�췡���˛����ջ�	%�c��!kw��R��^���.��eLi�x�&`��J-�vj��^�}��Ox@���4�
���lPs��.�nXMoN*�W�|������N����A�4ğkm ��.t�(�di��ƀ�������N(p��M$pN�:tT�Mi����Z}."���]�"���~%�L$c2�n۽�+v/ѷ�C���g��N�N>q�G�	�� n������t�ɸ����8�-�ݘ�ǳ$N}�\���Y����������k:(������N|�$g}o��\
.������|\���|)��Z�36�H�!�;�l�e�R�Xx��H:���eZ	�F��a`�K����x��ޝ�,����C��a�B�\Ji ���7��"-k]0�j�g�PհԂu��[#�s�D��TW����wP�Qk,��ee����k�k�`5���ɏs�+N�J�j�[n�.�~l���KY�=-t�
�'B=d�_ �C�U�}���u���ڕ����pa�#	�M����/H�r��8��;�)�%�Y��n�pQC3?�I�Xe���<X4���
m��8����q`C��/�X����<��i=༙`�;��٥\��Sy� p�F{w��^)��G�D=����΀�ϓ�_�+�q�]�q�J��ӄ���/Z�Vx
K����|O} ��,x�e����X��D؆9��7
]%�wuL�u�����%�S�b
��cS< vM^ +#E�Pw��DEY��DP�=\`1I�?���Lx8E��<��$�3�. �}��������;�o�`XW|��)}[B��?�Q�AJ,���5��A��	�	�']y���_u��Y��$i�r%�^g$J��Gk7V�)�..!���oN�m��J��Г+w�&[]^l{��M.	{�7[���ϻ�7E����@uY=����޶�z����͠n� ��z��?Ve�%�L�σ���vp��SB=7��;�+c����7���%�n�μ7���,D�����u��Z��M����2xZ��/�Se��[Ц��'�yw��ޒ9�@�yzp�����t��Y�+1�~�����د#��U|e�8�,���1��[�C����M{�p�q�ǘ{�i�wA��u��O�S���6����4h�\(�7��_���w��4^a����I��i
)�0�����o��"�A�+���1�+�6�N"`
%�8���v��baӨ'�:W0�Ӕ��S����)��1:Qr?i3�5�C���Mmמ�r��7�h�zR�z�;68
��t�ؽZuN�}	7űЙ�N�{{�ɍ���Ȭ�+�J��zq��ILx�v@<�}\�u�Ǧ�Bi��r犍�N\=-��0�/}������ԥ�'�ѝ���%V$t�/[h�������Z�d��l#���+i�w}���Ls+3�������HL��zK�e�5G"�e6�O7q��?&�Ѹ{TI�C�zq(+��j_����Q$
d�ag9�{_ g7d��WG$���uG,c��z_M��QߞذVzEÕFA�.�!��x�a�_�A�ꆍ�s�Mw�9�����v�x3WY_����滕��kN<q��]J4�aH#�������,��W�����?ʍ��Y3�q)K&�ζ~�W�/Ee?���(��"�{3��n�g���k�A����{U64��v���e�Q�r�&���3��x`�;A�вO�uǑ��%V��C���I?�I��S
�=�8��]�c�fv����}�c��E?����
�ڐ�e�N��p�v)���?)�4_L	��g��F�!���W2���m�gq�C8hڿ�B���f-��,z�vXk��8�G:��a6X� �_��4�]�rS��I��!&��Q��yh_�=jevE�T)�`��~m#�x��-��p�u/v��������5��rY|�cƶ���#����K�z�E���a)���W����;��I7�<	m3�v�|�2����|�,��g0����SLtβ�+f�9�.ȂZ����Ў ��'C�4�����qC�~��T��������s�����c9�g��n񩣏� b������M2���bi°!��M<[ɧ��Sþ�Y1{��4HP��f�^_�vuӗ�\`�! &mω�YCμDj�B��iy�GR�hޞ���(3?�e"~�JI��ʻ��X�g��`��)��H10AwR,�°���&p���07����ҜM����Qx��eu��K6X�F�9.-@FX���>,Ŧ\I�p3�ɐ��A��YN�Z��{�3�H I����
�`'��/����|��b~��F{�S�9d�ʩ��J��s�ϯ}��آV�~G�ƾ;Al&�)aW�ev0*�,D�F$:�7]���M�d#ҫ��
��ٙ����~�cM̰���H��g ��S� �	�����[)J�^��c���՜ά'íQ�H�5Ok�=��S��J.b5}���mr�bmB�<iZkj?�2v��[�J����h�O{a�{�s7w�f��c�*�SU/�"{��β߽9�=�]:���o?'���wt/&?9�����]�+��ι-�hU�Y*?�R��o�����M����Q {�����r[�� ]��E��LP�8t��Z�Ĉ���7�*������1�`l'�@1wK��{x8t�vR��5u9�B����,�
�?���t~����"���Zn��&KA�#ш��X��:®�P�����w^��9� {Q%�aOt�ڱ��eY��{���!+��#��t?ہA�*äDJL�p�o���?'%T���Z6au�Es;FC�!��ڌ���l�m�����>�y��u�+y}�ҡ3hW n���̳DX�aA�˝�PB�e��I��F����ǳD�0N�d "- �G ���W���|��n���Ƨߝ�|��D)�nR��dILj�DXё�M.1~�W��#��a�� �bK��D���g]�_*T��5^N�B�yh�� ��������mv>��%+��V�q�a�t�(?��*.�]v[O�w@�8_+�<eJ�9~�������.�Bjs��R�ﴱ��7-YS�����e���E�M�Y�O�꼞�-!:�/�J�N��`�?�쮲��
F�Gks�}}M���D��E]PXv���/N+a�B(YN��!8o!ZT�잚��;}e��i�Kfc=]a����{�f�;?Hd)**R��{Н�L���z>N�o�Wo�� *��wt7��o7��5�����F�LN�1PBrV�p��ou]��;
ք7* ���qru9>&�wt�pQ���R�g0Ԭ�
-�2�)x��dΫ��e�E��T]�C8��[s����R��\->�1�B�%�[H���t��[���3HB�-=��I�A�"�����6zl(����:t�n ��3����E���"�{BE%�J�P�
Vֵ�U�b�sկq)�eU�thF�
/��R����u/p���C(�������8�("Ɓ򳁄j��@����Q$�m�����xAVB��6/E�,3����.S�zno% D�\���Ё̜0zH��n��Ѩ�Bj�	��b�i	f4,3�pz�yۀ��
!��eb��|�Z��2wF��AB:����9�W���
Բ��l����[�b�z1�&|_C��*�ķsm�ٶAy�A6��`�~����xB��a,k4S5:����U���om���x;���lNJ�O ��6�g]ƒ5��4�8�l|��u�l�&̵ў&�oG����-�q�����{��ŧ�y��I�+�@�t����쉕&�ث�����[�,@�<�d�xYl���{st죮
[�x��W�Oâ9�h'�q6��V<���׽	����$
�̼1a�T?`���uŃ5��� -���n4�P�E��9�\��Qܻ��>�U�6ސF���;���kK3��Yr����q=����m����F��"�ZЪ�G�Q���`���%��0m�r��U�h}zr�\m=y�l�c��7��I
s�����?q�T�Ϧ�T�:@�1��	����{>�	��m��N���/�AV�Chm��!�_��uPA:�tMt ����iP^��Ҥ���R#�ȋ/�	n�ƸqGk�'�g�q�5��,�.��Qx{s����0A�&���+։MX���8���c����#V�
o#���u3F��/����B���݊������}ɍ_G�����h��zp�Ó�_���pK�h2dP�A�拆���L�f���o�՞�>.j2�!�Io��$8����f&���}p���=�%Қ���-�:���6��G��������a�;���Z�8T7\��KN�'��4�ťx{�0!yl�`�i?�H�ҧ+R��g�˅�lp�<���Z ���$�������^�9�*3ʫ��hg����)��DN��0�le�n��r�$�C�-�A��-a�(GQj���N)�!*���T��q��}t��X�j,Kˉ��j��
cq�R����4�ԝ�����;+��ˌO�v�����}>����NZ���y1tB�3�_%����*BUfo6�ʵx�n���қ�6�+#��I�_ �ճ��(}2f�:�?�w����_Zo.�^I*�N��Bɑ_�4u;y��cH��WF4�����Y\����>�p1�װ|qyo��:ѻ�j�o�%0�q	݁0��0E��X7<��=��u�cf�/���)�;�MY�Ӂ���#S��K�
uWP��Q�)�q�E˪���d�>�x,��\�Kq���؍�<NoRt�i{�9o�s@q��n��ؚ��R���T�ܷ�g�Ӭ��{��~���t����a1�1��"$�@ou���"j'4��V��p��Ό�	D�l���'��~��D���,���G4Wgi�p,ć��u�o\��߹�`rHs@��J�j�ն�M�Y��-,P�ۖ|��ь�Y��a�U�������&3S�f�p�dԂ|ò�~�B�aez9<�v���C$A^�k3��f��"NБ磾f���]ţ�rzҶ�Apv4���� 3��G����M�R���#w�IG���&��2�i�ś��W�UE�I���Y��x�$
x��z��!p�e7h�r�w�r�����,��g�H�A<������UX;	��Lf%����\����3�h�쐢z�)�]���ey9�1MRr�>Y��d7�P�vSq�<1�RR.MC%L�'3���K{ɇs'�b���ؠ���1Z��U��ϙ��曽���քG�z?��t�]sx{w�s��L<ޭ��U�O�h��i]�4��-�,	9�9��-up� "��g�s���z��>S�'}����r��� �ښ`R'k�G�xl.���/;�U�����
#��ZiO��?ǼO���k��������_����Z��Ђ�O/��{I=��nz*O����z
����ځ���uTybJ��8�~� ڝ��|�J�~#.Nq�;�q��ZtԭioӤ��A(����˩�¬�?�<dT��V�ŎՄ����vVۗ�;720��?5�R����\�楿�0D(w��ox�I�:���ٱ��jg�;�J����b��+R�j�/HR=ﮨ���e��(��*�~����xC�٣Sr5�	a��b3���'� �ki���#gx�j�(>+O݀s��W|$ �M jҤҿ&0��:�WvD���(�U�׭*��h�	�T�>Y{f^�]Y�~�2@OCU]�����s�Ћe��ў\��^�i괇���z��e��fj[�dњ;�a5�~'�����zv��"�S��Iw�a��P�����mI}�6�3I��j�ό���"�`����D�,
n)	�b�7�}s�4�ES�$!V�j�%��0֛�`H�"�������a��\U^��1�) �#��� >���l9�ޜ��� �Z�)��� ���ҝ��Q�WSA*M���S�De�qR�d�h�V�tU���;��g�����Q��%j~&vl��A`�d$cC0�� ������~縐	�5թKM�ť��"K5�{�V����v8h��l��j*�L=��W�X݁=�	B�Q����
)����x�y2�=<8�=����xq�ں�4u��b��ӱ��OZ��˗���8�V��ly���>�ou�|������0����O8�	��1��撇��S!�j�������W��4�R�<��=SYJq��<�c��,	e���y��.�i�JFy�k��?�s�&WW5��S�+5�V�Rp��1�'��2�[�>�˞�$��%LN�?F!���9������ �䈌�d�zB`I*D��J���n�|>��y+'��T��?�\6	���]�HYE��)>�\����ߛ�u[�_�:��x�B�t�b��aQ�����k��/-$�Wq���,	���;Tle�o����{Ο�P�]�շ� _��D	����@)��z�b��,�7�HK`�p�at_�z��ݽT�)/ѐY�Y��	�.k�:$��[F����l�i-�F�8���9y�Wq�}3컭CIr_�(��$2Z<=�o�Kc�x��M��\���CrA��?>`�C�.�K�匁b��s9��\��
�"������4Q��GBW�0�'� $�	��E#�縐]yC��x=�d�!�~�ڣ��y=���(k{ds4��)��ì!��ה&��E��:v�����`��i�#\|��@�T��%�u�B*W�^�t�����F:Ot�ϣؐ>����*�� �`)2��&?�V���<S#�dE��"��`g]��-=$�\�UI����]F���O�"�(Δr5�{6�!O�\�&��?�!��������6r!�cO����Z+qL�"u#���3N�k��f�6	U1�[0J��yy1�e��W�{_�ԥl�>N����;
�]�/�y�u䕶��S~㲢vo�t`N�i�9TnRW���� �[�Y��Q�b�7S�@���O]`#��6�C�3tbh,��q�9?~ �B��Y�^����]�Az�S�Q�8O��H%��tE�Σ��9oϟ��<gV_ԋ�ؓ��iTЎ��F������=e�\���/��V�����]QHU�+��s4�E�����v��0�a3��+�_VS#�N�־�]���_�dN��7#YI�a�\P]����ѷ��ߙ�	<Cy�7 \<�5�~�f7dF;TSH��H�|Ɓd���wN�u�'�/A%P�ߡ�H�;3��dP:SD�%8����Oq��g��~�e{M	���p�{
v7��k?k��DQ��yC�?��#�T=�3�j�H�7��s�j���3����0�Y���8��F��A��$%����n7�-D��Sc5�RCm��tl�g#v^�X���|7`���6��Ἓ]2ߐ}-rg����Q;�����m�b��ڎ�g��tZ�p�<a��YJ�wk%P�	��x���o��i�L�ŹKw�+��@]H���JX�;�;	�`58
�D J���"M�Yr�	�F��ޭn�@K-^����3�����ԧGp�VG�2ȬCumQ�&�cI�3� 'rUS;�d�U��f��:�#b�^4���K���"@��|��6^�S���s���/ 4�߬)� �12����O��
E8�����e�v�~1���@��S�FEz�F��+�i���щ��!"`��\G�p
f5�v?p�/v&_:57,��>��$���0�m��:��`p����� d����6:A+�#��I�Y6�v禒�SC7���Kh�� 4�$��,륂���9���&q�,1}n�i�)̪�o�ʉ i���N<�yR��/t*O�[���fƝ-��@��fL��!���*���(�Q�#�cg�T{@'�M��ct�l,�Zv�/�o����3d�n�9l��Y$��x�%n��#��U�A���q\�0���6��'�6��T1ۑ��+��r�.Y�s�M6�m�~"Vv,2UlY��>o�c�f��
��(�A�`\��;�H�@����^H���B|�S������il�ܷ���`�S��s��'�jjX���Z��&
,�:Ɇ>��~7�pΗv/E(��٧���N�#O���5���]P.O�ؑF��&��k�s0���g��-��<��G��<s���W���h��GK��l.m�%B�+A���e˚�t���}uC��,����]��"a4��7Ӊ����("�_m���.ⅇH�������#?��&s�;��88�F�)�!�Kz��4W�)֛>�Y�Rz�08+���1
�c���SM�|rD~��� A�&w�g��LҼ�֟,1h�7K񂟧:�\���j҄��ߚ�~���X��KX�`���U��
_��� ��+��t���A��Uz�%�岿|�y_
	ӳ�C�~{�-��uM���.?��\��xœ���5X�Z~�^CkZQM�eM��֖��g�@Ԓ+OeqЅ��跍��X�3���PsXd_��u�^�r�z]�.)��c��&�K��֢��nnq���
׸6�[`�ٗ�0%���A�w@���;�Xśh�2�X��[ࢭ���k�t����y�[�s��6O�\��� ��8ȏ����3}��Y� ha�`�2�`�����0iv{��X���1���OӸ=F����a oQ^'j��!= �^�iR����k�R�@��Y"O�;�w���/���Ң��0�n�q����6v��@{�IǓ�E�k�z�];�h�ߤ��l�xg|������V\A1�����O��I���_M�faY�' 3?2 >9ܢ��@����H"3���ֲ-���O
����st�4����U *-�3/.g'0%��-�3>ީ H]���b]�UD᪫g�I�l;��	P�Yw��f��e�\D[�^�F65v��+���W=?9�"{�m�����׺QV��~2o�������axG�#B���C�(�%$օ��`�QD�p;���/�\?%����2a�-��Wl�}�9c8U�u�dVD�K.��`�T�Š���kš���Tx��*G���:�@��qTv�2ߞ�@���k�SHi����	ƈK}�E2�ser��i
���o��ӊ��'�H�!Dq�����ʾ�+���k3zif��T�7�|j�Pzb�I��)^N�a�^��6�o��O*ʗ�Sâ�(�!;b�{D�8���� m�i�}d����N40�m1h^u�*���`h�0�-��(�
:lVX� f���$�p��=���I�[i��ϥȻe�ym���6 �XvȺ�./b�5c��n���#%7낡�-4�D��C���G�V�T�u��?i4�J�4�0��U�\ۗ�)����N���@��T��}%w18K~7� Q-V�C@�v��A�f+P��y�E[�S
�C�V��$�D�9�^0��	�g�4C�s��Pϕ.�v<���J��+Hn!C
�������~�0��\�^�W���x��g�nץ�-�vJ-rt�m$q~8ϲ�D����+1t��6���S��@0�a��#�s�ˉ��u�������iz)P:��_]���t]�bNJ�h��H���Z�yI��T����kXw��{?�r$
�/��Z�B��6%��jH/�i�/�"��;$����Gɕ��~
՞0��̭�o4A���N$�z����: ��dW`'y��z0��<b��ªC�K�O���5�~�-�Lh�;����ܩ��z �����G�6!*6)>UU����mS�y��G�����q�@����L`����Җba>�ü���:L9~ G�/Q�1�.?=��`��#l��rO��%p��08��#j�q��j�*G���AW�>N��)�)���0�("M�����k�}�Ґ�m3�[��9�Ou��.�q�X妚�f��(��vy�IO�z|G�@Q*�Q>�#o���6k3$|JL�r���ガƙ2ϓ�3x���"��)7��E��8�|&�p1��@��-�s��������0ma��T8��K�1O�+YC8�=��*�coʆO�sﳰ7CR�A�;6z�."�kn�;s�F�g %�Sf�=�3��)����fi��`�w���ӹ��P��2�J�p�cS�2Z}��Np
]l7��nf .mv��wd�P��d	*�E]�8���Zog����_f�ƘߘM���(��zU��3�����ܗ�'ux�ܼ��`׭�M�����d��	��[9!*��;@���t���mE���.$a_S�';Ԫ�ԫ���f�w@""����k��mFс�o�nެ��
.+/4@�v�1:�vj����_#�簎�u$uI�l�HQ0��j�\�MzX+�'� 	$�J��©��Y���m�K�%~��!Ф+sH��7=O�Ls"Ѻ"'�Aj/6fB,���>��y���Qk��tK���u) WJ�0��%����
#Dt�#J���˘�G�$��ڰ���QG^�S�%�g��[�_�}�'�+�Z�ǜQP4q9�C�U�.N�y)���ֽq�@ŭi��p�1 (���rqE�qq�^�,͎/��¯*F�=�\� ���T�Q�Ua�Mu�MvO���?����X�E���;|`@��6�Q�T�,_�����n�@����H��kUf�>>�0��-X�l�h+x_��	e�	l�Fշ)�o�숐1̔�/�����g�l;y"��B��ꗍ�5T.á�B�7��C�V>�FZ�&D�eg��C��?%_1�iM_z=a4�wE*��ɛ7���{1�(��&�~�V��M�㧃��`t��:	=��S���/��iJXg�9�{y+�5+�?�/���6;�t��aK��F����^�%t�	0�xK�/�� �I��&��+_vA��\Ƚ�}��g�M�6�a���'��4Gu�r�f�CԿ�-F�}9=~\Ǆ$�B<�m�	q���aZ�3�Ub�I%�������A������{�U_�{�|�u��bJ�����uR�r����g�I�S�M��\���T�>��b5Ɏ����㗕V��t<���)��2�rt��	⊟��߯Tj5�0�����,;�N֨�����$�!�����V0������
W��3I��8!��2~��)�#6y�qcq?8���)�h����#D���H\!p{ ߩ�., ��������� �"�X��a�5�����~!o��6r/��I'�T���3�ъ��kX�������v{6:�?�
*q�DIZ�ǐ%�wI���HP�H��ŀ����Qa>��Rm�J"F;�BձDڿ�ۋ
���� &�U��ȟ�9,��5]}0g��,�8tĞ�"0�6��׉-���������{T���:�gS z�sI��\SJPKc�D\&!�]�\�4;/�H�~��S��q[P�˱�WӤ�����	�m�8[��p�"���G� xg�+.d&R@�`m}v��L��ٖ�F�Ѵ�Y	��#���?��A�-��e��/[
h�[ ��8t�`�$̣AV"��YI��y���ė� /1D:����w{��Fu�>��$�CRT�U��K� ǧ��
w�7f`�J���8D�������%4�U����f<S��������Q;Bܪ���
3z��+��E�
D�E��#����	��l�[�63�K��N0x
6x�bV�bއ 	��Ú�����#�U��.˪H��>� �ܭ- ��q��q�Yv1<��,��_��uVP=�_�q��b�[�g,�j��(��m�lg&�%�WE����?�q�pUC(`�[�/��$������J#f:Ȁ�y�,d�Qm)!���H5�o��f婞���B�ެ�`�?~����|�����y��C?�@����ϼ�H��V#�_��Ä���=��h����+�CF����U�p[��G>dр���)/UdC��_iP��X��]�Qw�%!Ȩ�#��e�Ƶ����CG$�+z���'�V[^�F�1g3�HfJԲ�r_k�ޡ˯��6�vV!��WZ%��4�� ��b�8>e�0���C���Ȧ�B2s�L�An+�%��Cڅ0I�{Y59@U���� ^e�WS�?6L�%�2:L�}8��q{�k��{����i.�V�ލ
�mD8�T1���:�k�UH���OS���ƀ*�xO�f�83X�+�_a5_ե�br]{֝f�eF�yv*�֊����ۂD���椌XO��k�WB�5���>���f(:�w\6kh����R��$���T�<���-0�)_lZᑙ+��Ե^��I�М��t��:�s�7��c���O��8����!>, ��u�l�9�r��Z�90a��^Wl~4-X��4�u��N,��v ɗ��J�UƇ7��b�t�~�v+A�^�{ާ�V��-q���f퟇x��j�׿a
t��N���(2�0T��c`����=�6�N�pվ0�U�`�/a�
{�#P����njI9e�ݰ�i�9���I��&���z�FV.�>E�u�T�6��#�C�����P�� (3��V��B�Z����x��3k����σ��ɢO���p�ꬆ��a�[a���a�@��4�����9��+.�����Biik��J��l8YxÇ ?Zt�i��d�X��7��v�Ϧ�*��]=�����f�]���+XH�)Byl�A�u�4���$�0�I9��Co1�)�Ƨ�i���:N��,�7-a3FsBִ�*"��T~8�ل�ve�u�j��i��#.;,��N K�Z`��0�:�;�ՙ����z��(�'^!.��Y0gj(���E���*/��=밸0�[�,0?^��\|��C��5��gF��CG5�����{�P��� $s�L���A�}~x�(���y��U�F�7e- 
%w,lr|��k��v����<)�L����u7�����d��O�Y�Je)}-���<��,�}9�*ӉC�cţ]3�k�C}��+��A��3H�j��%�@�׬+k����J�S/�z	���/(���v`k&�_m�~\�����4U����ΠN�8�۱X�`S�	0VA�8��%y�<����H̲a�4��=� ��k�p<��E(1-�04�-i��>'`�#�(���e���|����I��\~m�6�Fg�x�-��r�E��Ӯ�p��f�y���ݮ�8p

�|�� ��VVr�y��j��e<���-<�B��x����j�b}�E0���xb��M
�t�[u@����W����4OH^�.� Ro�� ��i6����}C-J��K�d��%�JӎeD�C�DY�ֈ���aF~ +w������S��x0\�V��?P)he�E9�������aP��+\4�:�����Wx=�:/Ԉu9�s uOa;�a�v��e�V�V�I���Qml:���r� �&T�P�����ǧ>!eV�J,�E�J|��u�����u�����̕z��5{�/�*�]si;j�O	jU���Xy�$y�]��!>RΪ���4a̧+D���A�+

������sXÅ�� �H�t��e�Gi�N�c���_�I��jC���k�}[�X�^��f�}�'�r��Ƶ{���`��l���m-�N�
�#�Z��7��c�9?�Eh��s�g"�7U��X�I��d��WP��3M^�vkס<>�� ����BD���y�Z���uϐ�Q��oND�������!�R�[� �&��`QZs/uF2s�s��Fm�p|)�v	l��ƪ��
����E;*��򓕶D8�� zEXX\vJ�k�v���`.�ſe���~�*HJb���[�H�f��"���Oa��7��*d.i���e��܁|���)4D�p}=��0)4g��_>i��o��?�>(H�`���6�s��IhP�[u�7��a�`ե.{�JŸ��Cq 2�E��c�nc��w��.$�[Jٳ�[܀�뼯�����!K�P�#�b<��x6'Qs�����-�;�]���U7�٫&|�O�M�x<��B��#�pv��9.x����Vu�!(0����F;p`�꛸���%z=9?�{���+
�����~
��U��-pn�����k�S�����3/���o�b��Df�V%�q3�+�'����d#�ſ	�6��7o?��0���U����y7c�Y0�n�
ɲn���M�T[
ힰÿ������A�)�R`d�fв�!�V�D��B�o���200��+��jA�ы�nG�lT ]%����O�Dg<Bt/�_gO�$��r����)�~_�G~�QP�QG�_���5m�� �^��®U�ZNG��xs�m�w&NU5t���+F�MaL[�����vң���>�z�Cf��>`��:ǁ����~��]K"�|��iI���Li�L0�A�s��C�zV����h�s{݆������|(Y5���;y��T��-�^�c|�+�<O-c�i���򞗼m$�-x��,����`v|pY�$5�4!3�m�%����d�(��+�/�*��0 :i�ɖ� �{�ı3�S4����SCg ۻ �C����5�r� ���Qd��99'f��I���Aj��� H-4	w��E�E�I��$��H2�Hk<����㍳�K�u|�I�^n>�i��k5 6�RA��U���`d�ΥT k�)fC/:��8����j'�"����7��!&e�N9�SiRl۫�P6�F6���5ֿ�z�b��gd�3�/`4��P�+l�P��V�U\��gW�{�=a�����iZ�͊
���F]�D�m�ԛ�_Z���������J��z/f������+W���^\�f�ۡ,�̄�>G9Aoi>���v�{ӗ���p��y��Z�#����9fBo���w	4ޠ3��V9�%��_�l�����z�!�}:g��q�I2��/&"Z� �h��ږQҺo�GMZ�:�#�?��!�9�	pޚhi�a���z�b_5����S�mGK,��{�.�w#dQK��Si���6M^�x5�-��ݑ���z+ }�j����O�4^yQ9����ujձSʌ���$q�?��~�ar��ѥ��
�`ެG������yB�M`�?3���W~��[}�:�C�0�����pH�m=��ŀ�d���hI��l���2	������cA��#I�蕳����g3c��?���4UE�]��i�4�'9N�(��t��87�!ΐ�<�����_���j��Y�NIm��~�}E�.@�t|ͺܻW��,`������v$U]�b���>�:0Q3�
�T�;��!|X��ء�,_�_v����;<K��I��Ҥ6� 2��Nn����p�
THyD0�g�T-�0�\�}�S��A�i�Կm0ha��m.�e���^��L�Z�����P4��p�Kh�^�K�0ެ�f_�+��e����y���ѯ.b�վ��J�L��]E�t��z'����R�d]t6��6�F{��)�����+#4!>�wc�,��FJ��\�( zk�ބ��m�ƞf,a�eh8��	^�M[�\Ek�ҁ���\�(v��8R�F��F0�"���PQ��+KU���m
��|r�L0,�p�.C�z���χ���&E������5�L�[�z� Q,ҵW<��O��%aՌ�����$�R84��)7XT��:Z�}x�����G��	h��Ը��C�7�ӓ
��U<7E�.����K�5I%��׍ҫ�<Bأ}�
3���k������_f`b�S�����xU�p�ȃ�;�VX�=+��~?WN�R0�MJC�;�j�CJ�Xܒ�nv�"@��e���s����H��A^��b��=������9 lޘ`v��Z�����n0Xl��r.��AHx�p���&�{�p�<b6 f"���
���3�h�]&�{�3nG�wwP���U�e����%�"Kh�s��0�*���.o��.i�����Y��L�i�K���]���~���!�T��&d}�o<���N��!�@oA@�g گ
b���&1�}ϭ	�#R�4�6���2'�-)�kT��U����[T�xMh��cS��ay��e�p��w:ɮ�RN�uH�$e�z�ıǊ9
�vŵH�2iJ��A�s�Ր�������jྐ`�8��5ᥲ�IK����
�����|u4�/����TӐI!��#	`�q�;��B�:���=)u"�t�@���!`^�r:FXTf���Z�ti|Kᮈp1̧2�����TB�
P�<9�N�+O���P�K�#	������V�{x�ȱdI��R6QA�!R�7�R��C��γm�q��u�E���+��<�5�ּs�>�����)e���/xc��}E�"�OD&�lv�,:��GZN �P-�
>�����芰VXٓ�$x�������MN���2����}k�4}�,�n~���g��< �~CqN�0ʑ3�Q��� ̈́^?��Y&���|�yZYџR���1������B�a�b�>�Vz�q�$�����C�Wٹ�+�Ձ�f2�0�>+��@7�zLȶΎ^�g �oC�=]�GFi��p\d�Oo��'k��5��Ot��i%cg59���*~Z��?I��j���k��EaA�a6�""�d�!�~�[l�d)maw��F.���Ѷ��[-+���Կ6pKu�E�r���>�e�LՏT�z�7�`���]��t��河��1㾣e��H�yglc"·��w+�둢U�$6�J�܉EP6'#�:I;hhx TF'��]�D�6�O7Bj�"j�X<�J�75��\�M���+��%0�4�_]��qj�d}�_%B�L��H8���	�����$�F�$_��1E�tx{n����U�H���P �g^5���&��#F/5w;���8Z�����"������
ժKi���c���K�"2":�h���1��ڼ����%�U���c�j��҆z��Q?�j5�za"�"fR���v#�kܟ,��@��J���{�`�"�3@����p����ߨ$�K�qw��*�@u�Ǳ�����<��#��|tj�`k��2��Y����^j����[�2Ҁ�����,�D,]<����X�����?}2�xYB��*�0�O�C �lM(�\`��Ȅ�F0����vq#��wdF�_dT�\	��f�'��m�8;�U7�����.����(m嵞���:�'A	�g��fN#@�u	���P�ۊ� �� vi�vsA����N�� ��V�f����&"K���q��4�h8���Z����*�-�g�F:����[����̠��D�X�)u���,4J�\�����zϳtL�A�I�a�� Ơ�#Mw`hy���4��N�
�ʣКw^Tl�E�.Ӗ����7/$�Ib�i���R�V(�9�s,O�|����rn؏���.�N�����ȉŅ(�D��\��(��˦��ɔ^ fvR�|�m��'�n���px�I�S��Ww�RZ�����O��K`&9���
�?�Xu�Y� �Υ�!if�
���1<�irCF5�>�]�Yͩ��ctc�ʤ�0i�G� 倧� ���J��v���[�"��!B�K��UpJ�]/��9$e@4>ڜ�_�}�M�ڕ��"/v��̈́�s6�H�4��@��_���Bu5�s���fW��)_u��Ҡ=�n?���i{쏮�y?~�4p?���{�%E��$p"�u�c;ɎBO�2��8�	��k��D�byM��Շ[��Ĝn�*�V��,��]�y|.N�9��mv����S>�y-����j$q�r��,S�i3�t�Y��i�4.a�p~�/�x��p�y�?>�ߔ�8 z�jUpw|�t��Du^�]d}9�"��yl5OA�:��u����Z�$F�tFP~�� qJ��r�
$Y#�-X�7��>}<�X���^Qio�o���&���~�s��44ߙT��ғ���N�]���MMf��a�~.���k�(Ј�8T-��<���d��b*6*����}S9� D��I�P�(�\�r5��N8������k`X��֝ p����G�^��i�fMB�M���N�վ[��I��O��sEܤ-Ι�\�	V�\���G�,��ϘnO�<>��r>uHͼ�\�)�6ﲤ�c�^k�Jp��v����a��rlp��(AU����