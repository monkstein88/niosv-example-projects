��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���eULuC�`�g��?77�İ�4�u�K�̬z�7ٝ�O S�' �#ͮ�t5b�,4�#��<V�R��y�\�����|T�����s����V^�A��󅎽�D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a���]N��} ��ַ��ՀC�_
�j!�x�vF�AB����:!�Z��"_z��Ʒ��ԐY]V�n�����,3A���uN��m����'�/Pʒ;��:�"�ܼ@�GB��>�P�=(4�w�o\�
 �J�F����%Ɩ^x���v��X
�U�����%.>�2ڠ4x�ۗ49��Nx`hSTv,2�Zv��3�Hqn�;�K�O�X"ۨ���2M�C�J۟��	U0�!��|�vv�2��;�L�-������޸����2����_�w��:UU^�Fmݦ�+��EIp�-^O�f)�z�5\X��l:|�wǐXx�7 ��Y�)����	�v�	�w m}���΂C��m���{;�.|N����[�B55����=���N�ʭ���QdOZ1;���wN��f��{;��+�D%�^~ς���ve�Q��d�A���k�Ȋ�#�(���3C���
^P�a������B9�~8�+�Vc�|���W��U]�Ҡ������p?Z6/��ԤQ�ƀu�
l�	�����m�4�7�1���3 ��C�okDF%r(���Gu�_x-���eKw���G*�5���~~7�
$�%���ޚz�g����*�/ �'ƌ(�W�Ӵa5"�X��G
���W�=D�,�KOӧ�G=j���O���镸ɮ�Wܿڶ)�Q;��H~S2&J)�j{��+[���c5A�����nf�^�5���Ka�j~&H��Q`W ��E����=LbMr5v��i�S�ZK��]ɶzD���Vt��p���@�r?M˰���7��]l2}��s�Ķ	�`�����:�����h^]������ۼ�ĸ-2^d�������O�֚�8K���7BUdoPMTu{n1��(�j���O�?�wkֲ	+���Pk|�A�#늩�2��k��d�)��!�n�c���gy �����!B��_j�J�v�,=٭�)�j�OAkٲZtju5�|���f0����i펣BS�B�N2��W���8#{��Pe�
�Z��0�K��I�~��op��tu��m."#���t.I���c\V�����I�v��d��8�������\��:��.��)/���GC|�ñ{����$���/�Wkf���	�V��jv-����T��#��w߷�=�_4҆�og[R_<�<�Y��I
��b�՘�BjcdOW��-�;	�����&��KQC�7����g��h�(��{/�tli�+#5�3�듷d��<p�>>M����Ty5�Q?�wWBH&>A,
��C# ��+졜;@���U���y}��s��D��~Ct���9R׽8��؜���Vxٶ��0�1��=C��P���ˡ]��?�XP�ؾ��#m�8+n��Jf�(���'�(�:�˿��|A���n���"(�Qw$��w&�� �?�I�r���\�����@R._m�8B��R�[?�	�R`$���{$s��r�lU�ű��]k��d�u_ Ƀ4�絈3��Q�� vӓu@�(È�?��� j���:;ֺ�V�Ec_l=S���uX��Ma	�f�8N��y��g̻���㓷*{@Z�V�$���}u�>�ۄW�=�98�+��,�r�?bH2�R(]�QXE'�$�=Z��/��X��ݷU�O/J���or��sdѼ�<���l����?NeU�_G:gT����'p�b�(J74���=����9_�����.��B�����0&}�9������?�PL�H�E�h�7"��ݳ�2��ż:�EԱ?�"��|�~u"��'�o��7��<nx��{��s��οC�ng�&?��;Y-�w����1�C��k�����2�l��UA��ֶp��|��Ȍ���;Wɼ��ie=d<O@Q� ��k#��������"��e�P�%9h��d�٥ \�M��b��� �*S��Bm`:B���}����DP��oq�	���f�t��w,V�D�yfl�絧<}��� ��3 ͔�g�������&�K���ϕ]*(c���h�h���$�8kO<��&��!�{����8�)�v��*|�;���ef��f�g2�#{'0��T�)�ZLyt�&��r����Y����n�X���#�b]#\�J4�M .~�����gZk��i�&���g;�gv��!�,X�v�	�w���lw[����HlɁ�{s��4HQ���=a��z�iE�;T?�����t O'G	�`�[H'm��%��-K�"��/TZ���`5Y�|�p�����̵˄��n'vd���A���Ԝ�����k���y�Ι���˼:�~���u�9�-Ru+��w�{��.�g5���e~~�Iu�+���"`9X;H�MwL�sA������+M9��kyo^Ә����'[���.���j�@Ÿ�"��?jth�
ـ����D<~Ag�p��T��?�K���e�lr	�ɧb�̘�Q^��Ô3�-X��9�oDJ[�
�i"I8�TUĦ��A��/HLTo����ۯB*\뗵Է����D�0�7֘Q�d�C�o��Q�RP�?���]m��c%3|�����pS��Y'�|�ۺ_I>z��r2��UbN��Fm)�.	"��L�?���\���|'C�]ю3����A���e:I�ȷy�^>���E7�V�ᛣ��i��� �m$��m6�$�@�e�V<=�G��3M����LU3��w@+�\���#�3�%�Oڴe�k�,F+`�x�(W�	h-h��l������gu$� �+�7İ�j�Q��_������mA�F�`��$��e	䠑&���~o8�Z��k�����T�lU��Z�w�PŠk`�(R$�k�ٶ���~U��4����y�6�)@&d�1:��oV;	��ΐ̨<�	���y�ô�j�W�r8��,��>�$Dl�	 5�����pة_a��5�Nu��� ��a$��';W�v����2+I���v!;�E!��쿯$_�?�g�u�r���l�Yi�^�	�-
.-L�FN5��:ꪬ��Ў@�uX�Pw7[��Eʍ�{���y�ۋ�m����~d:�G=~m���`�Y��DB-y��S�Q�?L�$պ�?�CV�<�"�{����>5a�H:��5-LGH)�����aSŅ=��x���^p{���LKC��^}]/!���H�,p���ubN`@����G*����ZH���1�-����9��'�t�hV=<$��.�wY-A��^c�8��!��W?��aQHY�i,�/�.k���l���ث�Ĕ�f�I�R{AnQ[q/�?H�2$�O!SZ�%T�ra'>��{jw������}h�|�.����W]�U~]tÁ�\���N�-���L�t!���V�@G�z�����1��y�Ǝܗ�w�8�C�ȍI��˻J葨9�uW�(�l��B%�Kɣ&��i��.�u���7�l�1;����y]���C��%$�b2x��S-�� ]2͒h6�P�t���n�¸�}�-KYE���+Z�D�s��O�����{����}�3~}�Va�#��$�lY�_�����A�_?H�C]�m9��dĵd��Z%���o�׾�B�I�R�c�3���/]��t�^�}��~pd>��|��2���Zf��l6wx|�[3�vD��e�0��� <j"��ʽ\FV7yh��a�I}�� �k�8�L. �u	#m�Ch��U���S/���	���7��NZ!�����*R����E�i��q��IL7R`���	AG\QH��z�G��p�H�٪�sH'���V6}�'<]���iH�e��� �G!ooJ�h��ʱX�kr��~�L�� ����������iH��I���X�[\�Z���/�c<��=��M�n0dR ����{Qw��	֗��,��8SuM��c���GwLavč�Ӆݸ.`�ʯ�!�/�o��,f F�}2�E-RLU���Fc-ֿ�g��A�$�S�1� "�_OjF��gY�rp�����w��X��	��nJ
�i�i�>�āUm�瑺���H����n4Qu�j�A�^z�����4���*�gH�܁�~��g2d� �}�=݄i��v�_˹�(�P�Dn6�Q���&CJ3i�o9���w|{M���h��(�:�T1E�/�f���ю�P�R"��Q�;Ҷm��i��5��(�8����˭��L�Z��!���XKug�Ux�!�ة�~ �6���2$����ꂯӔ��3T�KC13��� z�|G9�;ޡ���ޚ<s�}$*�2��\D*^�s�,PE�!�$r��S�xG<���Gv9<��s4�-B��L��Z��D��[�բ��4��vg�O�C�:R�R}���n QX�6<��a�KMVzO��v���޸��&m1��F�,%��<��Vw�;���9��Fԟ�&g�#�P\,��Tt��~>2���e���7��=�\����M�D����~�^ZRh���I�?�g�}|Ab@�ݹ��sm	�1�����pB�/8fx���xS�q���c�9 Ua�����{���ۉm�%i���Hp5�/���
���2fDq�}+ؕ����O�Ab� 5�CYGT�|l/4z?I��72K���7���塤A��eK�5Ka�a�%Wn����@I���B�&��I�r(!�	�� 5)�Nǵ�d��ϑ����8��!+E��$��\Xc����U�ԙ�G<?�
P4�Eb�n�ڴ�FF����V?"���n�/���>p�?if
[H�ǖ#>�(%�����Pr���������%�J�9���m�|~s��$�D�g/�2�SY�1(͝��֑b	Q��)��'*o.~qc��:���b���v������s�b�T̴;z��x�r� cЊ9��>P�/��
7�{�(���g�˜��$b����2��"�-FU7m��blbMm`Gz��ő�ݿ�=R+�b5�Aj�O0����{���C��.Y��������
w��w�N���q�*N�����d�#��q���`�m��e������y	��[���W��(Sr�=^+�yۺ��MzhFz��\ݤ�p̀�Ĵ2l&��b�u�Vm}ш�����ԣ8�\t��8��I����2�ˁ��^Uyy54�,*%�N��Y�#2�.x�	��&&�������qx�1r�X.Q1_.}M�(��]�C���o9�5�t+rl����G�׌��.cZ�<Ř5�_��'J����.^6oU6�������a�����hM.>f*����גv��P=$�zq�=�rѾf��A""�$m}�<Sq;
9� �A����f��k/0�U�ׄt�������nس�T�ydfL*;��l3�p���z��!�)�7���k}R^Ta>�T(3�HV ���)����>�x�~��Q<)��۸�;�	M����#�l=C%�x�]r4z�8��&�@Y98:)����Y�ױ�����B� ���� �`�L�.鳝C�o��:kBkp���_��m�2�^[�E�K*SY�h�9�Z�P�B{yh�T={���`�?�5�U�*=��(`���6�͹�#��aЛ	,JXfhKgV����8XyA^��������o���esg/�'���P(���
{���s(�sz���=&"k�iP���������2��^�lU9���"�M\LD�Tq�{BjR���n'G4C���q��7�����8�|˫��q���hm~?^@?S\g_Q@�sh���w�;�2�Pa�;5B�M�E�:��	,6C�[� ��<�G�d
���,-�a��FR��q*�c���r��K����o����ƕ��Ol�2y�^&�B��z��,>-RA:���|�0�!���^�#cv�u?T�h�3�a��}��z7B~'�3v��a�=w��_F�0y�����R�O��/S�Z�=���+S7�m����M𕥉�5S�>{�Q]�}U�0C�u���_[4p�t��4Tl$�A��rA�agz�Z׉��5�Aj��T|yC;aLY���T��>�}ݵ4MYl|*%�LIʅ�׌�����ă��)
}@l�S#5*�:�B�������4Vϛ�P]Wsv�v��O`e:��rp��)3"��͐���Z��@ 3"���ֆ_`8����~Jn7KH=�z�y��#-V�a� ܶb���<?Z]��[p�X���M����Eq���0֘c0d`��1R�r�w0S�&�m�mƚm`ԘG̽�.X����^��S��ٮǀ`���]���b!�sˮ੠n��pDfU�Fn�,V.P��[�Jc:Qi�Jdk)���3��Itr�&�޺��kRO���cܗ�/ɼ<���R���z �~C3"�h�Ǵ���5��y�P�VS|Wl�S���Sg�U���&�,�5����T~�hա�J
��g~d_.4ޢ2tI�L6�|�p�y���������{E��m��>��������[�I�I��v��2}��*�s�h�L��L�B�ir,�%��Z�w�����0j&�շe������|z+ z��A�x�œ�3����o"�BXV��NK�د8�z����Ƹ�=��~a��')�+����������Z�H�c4L�Ec���n+�����t�+�˴���{����N`�n�%�2w����MXgZ�IM�T�������L���₍�=X�܄+����NF��G�yYp�Xw1�Y�{�s|�s9�����움Bi2���6�Bg��>����]�ǩj�x�,���ET\���(^�s��c�3��u= ��b0w��5F_!�.~=�� ��dz����67g��E�j�C�� Q�D11W���Ձ�ɰ��:�st�:�Z���Y����>T�Τ�蠄۷�9i��||��%]�|z(�3�-Ʈ�w��S��;�M.�����y@t�CJ�^2�T 5��+�oT�p��ԫ���lI%p?pt�
:;&�̫
��d4�i}�+�iȅ	F�dqb��g��i5��R�%��R�@5�ϦQ� �e�[��-�U���c�T��[��f��07V�ϲ�9-8�PQINǋ�h�Z��B=2����Ξ�ZY����S��P����?m?�|�N=�m�@\(e�V���DZ�ע�l�9���˾���?��9����J�v��P�� �8d�Lm]�Vo��=ܮ[G9[������SE�|�3L0���Ƨ'FByz~���ڛG�Y�p�A�D�(�ק��;��fG���E�tS�P�W:J矸ZW�6W������&�ZC��c2��E��2�H�[�	"�f�IY�yC���S�g�u#�j1%R�q���L?�(N���������U���C�^�s��3��1LB��f�T�C�Ȗ��&ä��&��*�{��r��,�e� fa��_[�Q����!޼YPp�˛]��Wߝ.�k�1��;��1�)������U��|�B^�"�S��l���A��)u�j�����F햶���IYe+��������Gy���R�a��ݒ��h�Z�j��X��ѧ3��Y�F̬� �@�`�Yp�<x�Y#�M�ټ�KJMHY?ǒI�C�Տ���F�?��p�t��6a�[����C�
�x��;��`	��;�E��	�s���>�;R����QB�qW��G�ׁ����]I��9��6�dѭ��0a�=�l
1bW� /��&&nʕt�`+s�D���2}���K&�@(� NSX�[�
[ʼi�k{�a���A�A<;�X�ir) 1��S(�@�(n�>D�1���cA�oܓ�3�w�����t�H�/��^W���x�������X�7`�Y�$Tn���2ky�9��_1??�u�c
�Ԉ���m؇�~��B�֩Ls�~Bv�h7��m	�CN!S�sZ���\J�T�L�jF�t�}$2X$���ׇp^��j�F�
�s�/x�(~c)Enl���Z�KC��`�3��f��Ay�W9o!�VT�ZL�[3Lb}Ձ��d��/��"P�t (,{�i��s8`��T�`�Ȼ��;i�(O$]�J� 5����CE�H�B��hz�$A�$ѓ�>�����S+ɶ?��Ep���	�F�.���h�e4Bh�n
�0�8����1/v�A0����w����OHJHz�5��!��2�yA�����f�L10��O*��f?��(���]c�\�π��X>���/��R+��������_OJ��Ϭc2O�Y{��A�b|��̄�,��j�R\H�>?a�#�Y�"���'<�"�b�ʎ��6��U�����E� �/���%��:�t�����u<� ����(@RR��j��x�Ym��N���������4��QД�50�j�q����( q���陫x^m������5H_�h������k��@��)�J���$NT��:آC~�D�x�0�h�R��J��,ѥ��)\:kf!�}�,^��Pc=I���<�(&�s�|�rq�h��99�i������w|�R[�t�μw7�ݐ�m�$�&sI����BHJ"H��d��h�R7W�V�>�ׅ�1͍�q��7�G�	�}�k�ئ��q�;|}3{�;�c�1ar���0��3׋��.�ب�N�%y��� a�ևT�v
v��`F���.	�l�v�*�9x���-/�¢�g��ѭ��p4�q@T�~x�N�l�����w�����*��r�]kH\ e�x��d<�"ŋ!]�$(�D�.�FT��a�[7aTCX�d�'n��/�m�7ڨ�\3RG��.i7q�#�Z`k���	ɨ�ދ&�5��z���{U���Ul�B�-�ߠ�A:���ɣ�jvd��@L��ۘ*O�1&G���9�B_�bڋf[$ܺ����yq,�ޑTm�h���ٶ���{/������r�Wޟ�hn���(�Ŀ$�=��îu��D��[�8qժ]�W�+�R��Ƶ"�V���ej�kX���9[��䦋������@Y����x˖qZ9"����������d|�J���ʆ���6�����+b�"}��GχM���A�����)���A�{���%��(.*&N4��^W.2�|$��'��EK���,�aum��،KRћ� l�):aP�wcyy�F�v�@����<"L���Kc��]��w�g>7�=�
��UX@tg���0X��Tu�\�.�)&_B0\C���7��x�[�l�߸���|�t˯�����R椝@�Do�6;��I6@����ɹ�_�Hu�| ^^(�G�%��1���WBn�P^�h�-�%�O��3��u��@̩�5��n
3mZ
��o�חv؂}j����ڒn�q���|F�D�M?aB�u��M�(��2�|��Z�f��|%s��(��Us<�[2��.�{��_?i�ܾ!Jې|�}j�,�Z+X\��_ca��"�jR��N8�z�dEk�A��g~���S����Z
f��J�V�7�Dq��$=0<��3S9_�������Gm�ƱP��T[�� T��ER�+[�h~p�}�f�# ū��^�Bz��Bg�5&�\$�B�o͏�����<�o�I�F'b��`;`4z�ـc7ȫɽ��{�a�̸G�(�j���1��>��[������>��g>mSJo���/�AS�-��nGþ���7��f���E�ӳiVb^��
~ݼ������I�s萩,�S5������t���
S��捹�}�lD�ǊܰNy$X6���ɮBd�:�<�2��^���W?b�Ve�g�����_�%Y��׸km���~<�$��؍`tOb��4.��-�����áe���R��n�@���, 9�Ԡ+�lCM�T�������4Q	�%�V C��\�J4���8:�<�h��ө*K��^�[�hKJ�!���a�Q[��!����ut������tz��.Z�E8�E�[���T����^�B�n�͞��T��Z��~tf����k�MW҈L n���̘񉈯��p
إ��'���;�O�q%t�ZC�(\~KH&�Y����|9���w�^ޡ�aˣ%;�%Ƹ�����I�>�<�;�3
8L�5+�]�y����DĦ}���>�MO�jd~H��7g30�Q�2����ո22h������h�ʓ8�����Q����<��I��<��Ż��Hm���J����Ug-r�T��ub���rp��{#�
f���x-��;��!�z��&�uMG�tr;&�^��;�����_���`3�/Б ��C(N&�~銼//ɮ���C�=��i��MW�*<�{.XgQ����#��ժ�~zd;e��#�-<����"�X<����q2(whk5c�P���A��̂�������e�-��ʃT��]P�NbA$�4ܵtku�T�N;�
Ę��B(rҁ�%��0K�>Qaϒ��`I~cj˛ƯS�D�7x�4	8�D�ʣ�i��?�D�q�.���z\]D��8�������eXz���yR�1��(�Zz��\�A2&]+��&G� �ʍ�*{����cIH�����qO���ͱj=��T&���wG���J�2������K[�8~������#��ߚ�f��1ߎb��	��X̶�ޛ�i8����fQ]�G�������x���3���Cz�L�ړ�̟���LJ�뀢�$(-dU;s�z���(�#���津��l�JL����O�x-%��{˲��|��ZI�̶��x��|�-h#� r�3ý��0�;ڱ��PL�x�[��E0h�]n�7�J��haO�
��-ln���.5@�R"��p���V�sY�Z�w攖ֻ��@�x��O!}�;D:;���v��L�k[���F7ѐ��ID&e�U��a������tN�1��EQS�ۆa
�1I�:��)�c:��->�Z�ܳo�e���MykS�e�� A��*�<�菉-�WV�F�Š� L󞺹|��=Άy7l*�t��oYo��	P�W0�)0��x����RK���}2l�<}��_�v�h�/�%�-�u���*��;�@���{.��D�vҼ��1�M �~/	�P��Rt
��o�DA�|jE��ƣԇO�)�>?���H&%G����5�u�ݗ-{>��[w��~�o�ں3��un�y��c�K(&4U��e�������>p��~��d�=���	i�LI����ݒL$�ŀM�Ls}�Q��֞d�ɭrY�)���e��Q2GxK[ƎݯRD�0C%HQ����d&�}�q|@�_	����[������9:��s$�~2��S&��`�G��O�4�(���| F��N�<����$�mgC._Sf̝��_�N�,UAP�$�l�Řfȑ]�Zu{'�,�ouHa��m��5��v:�!@�_+�}a�0�a�絮g��6!(�$t�)�z2=�,����u�	hb6&A��Do!K�޸��,M�Oi�qXD�/Q���)&��H����fM��}HUpL����jeU�2G��?�v�O�fj�4��ˬ_S@e��q0��o��9\B�{篛fs�#0M�W�S��ϟ��D?h?�yfGr(�K�;��3I5��}�4�-��uSxqZC���U5��h9u��`Ϣ�4�Buʈ�f!��i�&x��2���g��e�PAVz
aiI�&v�B���wJ�)}��v�bt��@|�
7���-R{�-�k���k��x�(�*������Q��z���ox%~��{�\WE���߱]r8.��.f�j�rnJ]�D<D :��.��rZ\�\�����I
�^tŘ�6Z�1ݘ��,tw�<�r�Ĕ��}���!ky[�-D�*k�wh�o�D`�X�B�?} �:�K� <��_��V�2,[�Ct�.��s|��x�+(>����״�����B ������vR-�&5���b��2��� n�����=T�o$u���	A�3iw׃$Mߒ�C��0�ߡZ1�}���PNF���O��.S��eg~\3Z�H�f<dyO_�+���A�ކ��Gx4�c�us��N؅�"�'�"d���+����}�:u2��%r�χ�M	%�A�N4V��.@��]����@���T
��l		�P	��;�8��f��k��&ð(�������W�n�����Ƀ�N���R�^?�(qn(�6k)��h�
=&m_��P�ɦ�c{�(��NQJ=e�(:L�ĂݧU������T�U���$�Qq�䖘1��1��k"ă^�MK<pI�>]ZE?�=�Ua���D�K�l�����`c+a���_���|`j�������E̕ ��<b+m{.1`u���]�� ��U��w�b.�����ҩ���,��C��<K1.��s�xsozJ����l1�~�VN����S	�����o�0�c1G6O�oE��[�v=&;x�y�q�O�8¤`���M�1Fy7�:�'(T����5EM�S�����k�	'�{񚣁4�<��������^.�
#�H�<�������+�K)�.�=hg���p/Ť�J2n�0��PJ͵fh8�p��i����1�Y�-dm�8�c~ �dx3�+m+Yd��no9P����q�*OMȠY�����J?��@�� ��$!n������ 8�B�]���=H����̅�Uѐ�d�F�K�kp�0s�(�62y|��>%�3_����vM.��/�iX�"�.�\�Y
UPf}���vj�y�w�H��i]4��'��Xz3�;W��m+�\F<eƨH�9^f��s��@^ջG�H��3w�<�~�J�J��#�7�ݣ3ȝ���ڤ�R�7g) 9����'Og��m���=MQ	ɞ�����f્��7e�@�Wqױd�N9�c3R�w��=3Mr�	pm%�	����kL�f�y�s��̣�標�g�Uh$�����:�2��I�Baђ��������ܦx��p�g�g�Ӿ���8���?xώ�I�R�(�h�+�{&�v��K�Ոk���=�u�G�0�#�'B�n�*%�s�0o�zY�=H�߮��t@Yb��J:�\��B'����~�%c�V镻ԃ#��G	��hZ	j�cx&x��~}^$�������2��\Q�jd ��8���w9J�5�o_ғ����zp3|�:ґ��<Z�i�k�RS��tM�K]a��Z�J�J1:�w�!�-�:B`�oא
20�x���R�J�Q�	j
�Zw�v�G�g�b-00\68��������K	����W�A��"r�e�R7�1j�o| �j~���I=�P�/C���c�*^�i[�pk��ͤծw���u:�Jv���>���U}d������a<Oܹ�riQBuW�O�� �[:��"�d��TRn8�W��5~=>��M(ZR�����H���Kr�z�:�7�{n_o:���s���d���s{*�teG���(����j��UJ���0�cܮ��-�S��U4o֔����c�pFp���;f�c+OzN����4r���w�I��$8�������8���Q�6b�3��f�̛��b�&t�^�j����y&��75�<��������b��@��j;%�6��|ň[܈���y�#���,Y��Ns�rȥ��hj����
�j���'�r�+�dR�m���|�yrFB����a ���*җ�5�Ɇ�����&�����s��P�R$��c�=���;�1S6�%�����	�Ɔ���j����xP�=��1�J�x5�#�mv8]��-A��)����⣺j��m�Ԅ?�S���Eg�2m�Qj�Aq�W��ě��)���;�1���f;� ����gޫ�Y&���,�?��X8�XqC��/�;OG�e��H߈9!�?�*��m՘��+����c9��%����oa��()"0�"����˚�mh�@%Nl���AZ��;�0ʧ�Ι"7��X'�jp��b�e��2�\t{�³���z�{�������7-�6�3l��rI�݉$���9�P�z,�N�'�6�>���Ӷ7fe���$� ��<3 U��[�"�ܻ6�u��c��'��������&����=/i]Wܼ���k3�ˠuż&!�B,c�h�s�U�H.btx���q�c�`M	P�C>C?�ۣӡIo@I��R�7����?���\ �5>Ԧ�Ih��