��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���-ײ`�>��썅��NX�6�h�@.C��(n)�dm���R^%��ĵ0A��b�����D�i��������O?JS����ny�O���ͬ��󧻚�RE�g�:�c�$��^��)H}oѩ��R{�w�K@v�8"�~������ ��	'o'/@={�Iy�a��Q�y�'��UY�?�:���5^��F��2+�;VlV�ǦaR��"$R����".Wb7�C|V���:΋�p]����;r`�MNa����m�a�q��(rt5���us�*Q��<.���]m�3�nQ/,'d!���r��b�#���\�nA�X@��9Zg"��_�Kz��(Ho!r�[�6�JnK$3!�)�Iy��$�>��GՀ�Lm��uU)�j��Wd������Fׅg魱�������3]yE�h�'="�;���,�G�vQ����I�q�Vv�wٰ%wor����F �"ڇ:�+\��/[{ge��) 2��%Z���|�};����L����8��W�H0��..A�t�U?����B��&��&2���S�G'c1���2s�u�����<HI^įA�E�f)�����r�Ï<lfѽ��_�~j��R��]+�����L��%�w��JQp����d��_y~Θ���F�/��0-a?��?Q	jmO8�F��{Ƴ���W�[�ߧ�`RX�V�v04�����$Y�����Ĥ�2:jN�CcCH����}�F����ӌ&q��>�����G3�j+�jf���/,���ʙ�X���c_j��~�8�V�^z'�\�NP����VCa؋ۅ��`�dx����a��M5�T^�A} �l�)������4�Qaj�� �vb���d>��!��&Td�[�;�3������J��0Vo/*�n�,��8�T:b����a�Uh�!��׷u��T,�S�x��E�v	Z�)�6��xB��&g�+��G�}��l�Ѷ�i���s�u�x���.�����ω=�s��ϧ5�,<oC�iJ�/'��PԮU����`QsDu4�ic_̶�[feg������> ���7������ S��z�8��2
"���O�ӣ���aV�$[��Ez7��z6Kkxp�/�}��g�J�SΉc�E~J�g��a3�+��v���٤��V�w�=�q��)��jp=n|�L�c2��O1eba:- B�:T�3�K���X�|?�1�?�\�m�*�E�̂AA�iU�}�!ݞ�:1Ȥ�G���4��S
�T��Bb55AG%����R{y\�3��ݤw+8�L�H����
H�������5�&����=k��"�4�X�[�w<Se�3�0����A�z�H���)&�I��I*.2��&m�X�Y,祱	�cHs7�6�|�5��:���{Gŗ:u}�|�8Tt�0��E��`Q������C��#�?ŉФ��F�]�B���]�ɓ&��4�ye12-|�vo0��ՍLuaZb��FvH�Î� v���r��A�e2�(����i�H&D"�r猳K�~�sU�T�#�p�vU�ey��HMK�7�;���޻is�\���t+�����g���=Ҿ�w�\��=j��nAdRa_��G>��4_S6c�z�9l�{��I�T7�D)��~����e�P��9<S�b�:�{��w��`�~��1���al,[!���@	2yL�p�|��u��#���vGüX����qHgI}�����@�(縱&g*�����'u���Ь�D���B`_ɞ��pT�![��b��>�(W�P������(ޓzC\���l-8�p�lE3�3���4%���du�b~o�~�J �3��9��w6����Eu���3HT²yS������A-�4���O����������vDT�i�eݞ���y�[��l8�hoԗ�k}7��ׯ�j},e������v��-b!T>�DD'b˞#��#o�P���Wّ���(
�R�7>D�8����5��Z�R�Ǩh+�Q��fag�9�6����W��Gau"[TwЇx7��,ʻ4����C�kz(���'
wF��$�n4��ȁ�	
s�2���{��kL6����ȇ!��ɑ��}��5A٭my�#�+��R9�
iӒ�(��1x�^S*
8ށ,���LrL6�ɽ�	�&�ߥ��a�+&�7�P��r��dV"�bj��UԀ�9�-8<����i�Q��M=���:м�T'�$�-��b����2FW�:M�BE���� j����.�Y����h5���B�� K�ξ�V�� ���6��k���;�c4/��v�!��b�����d�F���kr��U{
����#����0�=^���	u�;�aH�^�0�V��5\