// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
pwK+lhLgZwg0A0jPs/5zhM+W3R7QbGujtlKHaEgXRqULqx4b+9FSDX0hW1ynCNVMRzaXORfyfN+o
jnq7rUa291jOQcR9pNDu7zgjz/AzQfQ18uh8r5vFxfDUChmI5bFNtI62s3v8SxYfKb4aL9/G6p4j
t2BKP7wI9NY8Wr55/JLZGXsrVHxKGgY8ISV6fbIZepR1VhIO3YFLvOfNieO4fff6b6o5GGcVkuMO
6SVG72j42nAlGJFoYlbxKfgN2oDjzFEQAPl3dAo5Ul57owR4fhc+w3esMvAUQrGGRYyIcmUd3VWZ
CgZiCskOTaxe0lxcp57BndvG77hGJMe+HRM/cg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3840)
uuHFdXNG+COs+UaQo7w+H8Ah/4bhZv8WAdra4HNxNR8Q6tAZKtIHimMqrkDwfoxMDr8NKhNYl4Hm
ploSSNwdFHe/MAHhH0UgW+0+cOBm2gNfMOfPrUpqb8s0xj56JpPojZpWKTgghqMa6ycskt5P33tk
blo2WLXjSrIMy5uq6EfTqjnjzXJulguyOTKFKeaWAyaUc9mDNUdfVc86C2M3BlJSKgc38csnp3np
EUdyZuLKFv6W/glThK1k0oGOSkUWGR4Tyu41rcDcDKo6gbu112g8EIwTkODhzAz4jMrmsyUJU7rf
dvrXs91/aQsZkW3KeTJeTzr543oHlJSLN67A7X/1QQsWZTwOQug9VeRc8cGOsjq2USPGMSz50hP1
xlgcys0ia46fMvDunoYS4saYlUft+HLwBDCpO8tzPcjKFBWo5zavfCKKRsnx+pM7uD9G9hBb87en
yfKcPl8oh/M3o3h8qzbbe8DHruwKtpf4IRe8rbrdvrKZggVa29ndI7UJYZWzNiwp1ZW/uf0EAjKJ
McIi+aSijRthdM2n01xqbZzmwdyWs6C8Kaukkq98HKu4iCU4BaS70IfRKvLk9hKoK/0xk0zTrPjv
AhDnRvCklMhIu9Vwp0wquXEpeyfSgonrHNgp0s1eRFRgbSQNqPyxzd8g80S+0/4xlckwmELTY4CL
D+AJC1D1brcQOqF+pu8SACdmOiymLAtS0tk38BxCMgFhJ6Ve4Hnuq/haIvG6bKJKxv2DshhIeNal
vHBJXPbE7fKLuEzs6PuBpXXNQ2Mvybwe0BuBTKfHEuPQSVB3+NVoaragChI3mNFuUFPncSTGYQlG
XRaX9h47r9iIWN0uES7UqQtwiCw11kcE2deGH/kffkHGeBTGslgu9VJQH+rvslG3xAhjyszGU4Hx
wM0gWUtpYXhdd+tpOBxwdKNh7Lcp0CwsicQrXQ/slqHydhJMTPj93a3s/zOOhns16JKpdVBd1riP
Z7IBQUKkdIQt1z3Z1K52jIUJyokzj7r8fqvz9bo+U3+3TMR+xldn4V2MCkT73qow7Zv3B3s7gsjt
RhvPo/Ih2p1OftqkLPyEu36ycdFTzTvwrxGX0Bk4KcSWWP1yhuy0d3nXQIaXNMYZsu7fovZSeDjR
LXMUFlpFSP95XLrZ9y+acSfPR9zFKY8k9TOB72e2nJqZPvBxyrIpEIsaedmeIGMgm2r5I8lORqYb
oDhFPtMOJzVL14MHPW5DUzYx4xjrrwoANpsBHISTt+F2u03KUfJDHq5jiVXZ3HX0MsuFCIT3u4VJ
9m225wJPa1BV5W/14YSAR6do7gCi6Z/xuIPG+V3UERwZoMKyeGQfxSm57iA/XYDEDzJLnef2Qu6J
ykFZnAqOz1B7rFYA/2YqYommnj18U1pK7Dto9BXRDpY+ir2VVC9i/8G5mtwzP7SLPSvSf5zd/iL0
jhNOMiY4EdpLq0BUH/Yj2xRO5LHiRL6/qSasa6tEWM7hQgTsEwySTkkV5JoKpBzvS+ljPndTqRnF
Yn19L9XywZqj/lrolpnHiuZozJHfO5GL5T9QlU/lWGyfyztW7WH7sIkPtqoBoCQA7Q5hcdeVh5FW
6Q6YqfAlJbbgImSbIVW0vifeRTuqOi9xDWeNVBxzo/iWptPymMGGV62ERI7KO4WTevmrEN99qn/v
g2QjeTJr5Ng7m+Y57s+bKfqF/wGRnk869ZYTPh26My+cql78CWh4M9Y+J+a62PyqzS5KzeyYVzK5
H5BPw1i//4TUqBqDCNRqbFMqn7c7aGX4IP+qU7VIJiTY0NPcZnmO7kjMGVWC58eiFAtQiGftj3cS
Q2SU6WEnOpZOHxwnAWDQXtg3uneCxFXLu1bp1/rVCqvRipW4b9eMitLi0ZHlG0Fotkl0moIhsdv9
Cqo+L3h6Gm+pBXpn6fHIYre6DyQ0yJe4o6eU4vMAVxMK4xo4n6BSVffoUWntmCUiI75jU+Erh8DD
vynSEojnOMfnfArbbGSXfTdfeENVdBNCTINcWjUe/macx05VqbBTuTIDv2SM0vzBVzmrN7EuIXK6
jx3SYEKNThY5mBskf0sMA6j3NFL+vrh+r0gEIUy9I0vaFddS/COdyjiO7MQ8kyI24/8HEedHzR+m
vBNMRBd5VBOn2nXhb97Yw2reblX+VFzmcq5Z53QTQNFCCo2lfN1o92VjDeoZ0mQ6PDYqxDO/jZT4
wOuTHmwLeg4gmYttKp1HYTRKCxOHehL5hqF4lIG+yqW28a0XSMHqT2wxkh7WMuMXq35ilEX5n4Pk
GnANSnIg4Cvr6ZK6OpB0hRtoWwy4QUyPLGyMh3nesLxhZtsaniImhtjX5VitiIxB5zTMW7vCRS28
70RKs4WU0KO0/vj4aq2C+YNh3sAWIaDGRzxaAk7f2iAnVJ8oMFRxMVNrCY1ysAVxL+3gWXEYBdhc
5koKrc5tkp5TxnM/5/gBfK2o0lUvS60rE/PPR9vLQ+MgyuVQG4ZD/18hI16b7fiQzST5s6wTp8kG
TKCJ0Zqgi9JrBLb7k9Anm+p1R9xM9x2GSEoPpVpDd6m+Qx1fy5QSM4FM4zIpWwoOuziqfF2RvYFs
hbRg0yXgAVkXqLhOiD8o2/M4ozM7/tHbzgO8PPF+tn1/2woqoQLD/svxsoaeIbdU3NAU2R6/guBB
66ezIPLso5f7lpXsQ52D597gQxrtF9agqujbRBrIVsmgeSXTYsWBpMx1PwTPdUZp2Zv/tBM+QXKX
Bj3exG7Pfm9iI8bMTaFHK89Gto1o/6UqrP1EoXnzxx9rmNDoIVduZQoalwF7zeZRCCfl73POP5fv
wBPefzAkxHmTbw2xk1l3M9DfPzZ22l851dPT/bIx4I73tiE9U1c0UsGqjKwDg4WuPr4fNTvQ8J7t
z9Kvfega4e4WYZz859KTLtY78phaF+XkiEI5G8vObCLD1Vy2rooCMgJRlVnf8YPhgokw/hoOwFnE
bcA4FQzClHPKtxsYfNj9QEMxVYAIWyrYC+Vi9iZ75FubEfogPfPMyKzCK+tjbJkWI9omZNX4FHL9
Sfl4ohBnroH+QMV3cT/KbC2Ocsn1E84XmQPlunTE10Kkgs1sC5YBFNoxk4dhbIL9j7U/vHSurDYs
t5OyaZ2KEsCltVFhbe0N85cZ5SoVwYC9RyJAjxga7o4lUENZv5Bfas6BHwu3ki1nJ1tr9MAZI1+N
xtyYtr3ZzH9k7FrtnS2ERzHsoMYqDjrRgKyyooZ2NkKDlM4v4E0r8Abnen+4bA9ArTu3lH6FHMYQ
HOGqt0Ha2tb3efrggixBXdurdBH99yKVqQp0Fsq21zT96JAIfcEwo21AjgHq1iJqkKEMvX6GDH+G
2urXVzRhkzFVOsiMyOgU9drUlCzO33TDLRr2NgTvyYtgSQW/2zqy0KSv2FjzkiyvCErkCKcsTUfU
lDj2MxpN9Cj1T+91YB5pn+JPVucA35HVC1BMjX3LDZcTHqsKAskWYj1QarcTlSVAkiUOvYo95JRG
q5FfbKQ3U9oVdVTQ7PQSCT5bJNP+aJEdgrk01Lvg6pu7h+akkfX1bluGsACFjjut1jMSgjPlTEVD
9ejtcgLwzJfDj4jsG3CDSh8GMjIImRt2ZWTUpZSkGEIT7/YFaKGhClgIsJDxMSgOzUj4uWezg7rl
qBBf5ZpUQDQvjrGsnnaHqsgFkzbQJ0sEBWXvLxMPS3a1v00S9j/zMa4mD+bMhJUzyB5IBmFFvmJF
NKWnBQxQzLvy27joIjWR7fd+hws8KM2tVQtdWh14DKGcMweeujFNJRrKzKyWkakj8otZ7KjnN2uc
ejZwQEcDy1hnyN+UpuF4nqS6dElO1uQUy7NoTjlPLDC2V7cg3G+c7VsjqG/EmT/W1+kW95ozTboe
wSkmo+0XdSILDfHz3Jr48vAdgEvF4VvdKn8P49/ZSSj6lhJebfk1EVNw6yildijEamNTBeiztY3y
2PQBjVhOWiC6jTMLYgcdi3QzB5A45i23heq5O5u7GxkFSfZ6HITO52IxdLYOq83PekYFDA6PlZrq
78LPNGrsa+Q0frLLbz9BIRxayHI3Cvs8Obq245jHOJRu6SH9O/sh+AN+EORtKGpQb8KMow8gbZq0
qEMnWyozyR9WnUyxlyahDnv1u72fLo1rXOBYGwfYXz0nds/1EqXGqAE9bzeN6pTuyWaXqUG4Gd3h
IGZXToEbsdtv8gQ7bFT3hGnhPTy9Wh7IXkwUswqzAb2CBHbVOVlNLX8dEe/SHaLrIRDA9dmgkJVe
YN0Z9lhTcWuwNLfnetuMh5/hxqSKSvEZDRhm3aWXQ/vxJ66Q39dm7DH3DTRYdoq3PbFb93iqlLTA
s+CsW2Qk8FRlOo7BTH6pQiPt+J//q+G91Bhy5udG9j4H0F8/DldDhmEKaPDspaBE+B3r/2q4Dy5M
Xz8aq37U27EhUFDUwKU7JUVDW2QD3batyCZ+7mK7m129zjglygbdZMfZuU24+mBByejBjcU1G683
55cU/Y4NWAXHhLuVxnn0wpSN3IxRL/aZ5l55x/HbOENSRMg9JL+Qw0q93EbLK7Vg2ooOGHhFXbqn
+HZksDeVkwNqbVbVkkixc8goVF3d8b7YXIPFwDZx56MB0WqE5x1qaEtBeAFt+I0NTH9eRAjYonUg
LnhjMskBBY1wyc5iKzhydh/SlB0kWLfHZVxxJGCn5g2laklGQwQdQ2jS1b4BG4vb1GVvFrkSGGRs
4A7QMZcGmIeO2qey0m6veYbd6wIb6gZMvg2Hj/gGX35WNUwkN4DA3cwZGRS2s17IV1o+ud4hFW6c
zQicQMHmjNMuW7tnSV27MMErEXcnr59DR4TV6s6Vz4q/fLvhWalqcqdqItir4IEMrXzKxJqKK29u
G9iDYpPhM8+FzKCn/L+XLAgufx0Z5fFC51OaqoZQbOubjxHvkOY1B24D81V9F6zZ06884h1d1l41
+19CRrJKJgOkxc+K1jjsawAPRuMVU1EYLsD+I1PzZ8ohh0r5tWrQrQxVNHgnqENR3z0EnnuoaXGZ
e6g8V8XRknHQ1RxSBiPoJj7bHo8XevW1bCv7rLUF2Yj8M2eKvb33PBQgGo+lVIyR7QYhnJOlLp17
JDuBPdVhVvV8PYnfBD89iN4kNUmS
`pragma protect end_protected
