// NIOSV_SOC.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module NIOSV_SOC (
		input  wire        altpll_clks_areset_in_export,            //               altpll_clks_areset_in.export
		output wire        altpll_clks_locked_out_export,           //              altpll_clks_locked_out.export
		output wire        altpll_clks_sdram_clk_clk,               //               altpll_clks_sdram_clk.clk
		output wire [12:0] ext_sdram_progmem_wire_addr,             //              ext_sdram_progmem_wire.addr
		output wire [1:0]  ext_sdram_progmem_wire_ba,               //                                    .ba
		output wire        ext_sdram_progmem_wire_cas_n,            //                                    .cas_n
		output wire        ext_sdram_progmem_wire_cke,              //                                    .cke
		output wire        ext_sdram_progmem_wire_cs_n,             //                                    .cs_n
		inout  wire [15:0] ext_sdram_progmem_wire_dq,               //                                    .dq
		output wire [1:0]  ext_sdram_progmem_wire_dqm,              //                                    .dqm
		output wire        ext_sdram_progmem_wire_ras_n,            //                                    .ras_n
		output wire        ext_sdram_progmem_wire_we_n,             //                                    .we_n
		input  wire        gpi0_butn_external_connection_export,    //       gpi0_butn_external_connection.export
		input  wire [3:0]  gpi1_dipsw_external_connection_export,   //      gpi1_dipsw_external_connection.export
		output wire [7:0]  gpo2_ledg_external_connection_export,    //       gpo2_ledg_external_connection.export
		input  wire        in_clock_bridge_clk_clk,                 //                 in_clock_bridge_clk.clk
		input  wire        in_reset_bridge_reset_reset_n,           //               in_reset_bridge_reset.reset_n
		input  wire        uart_serial_com_external_connection_rxd, // uart_serial_com_external_connection.rxd
		output wire        uart_serial_com_external_connection_txd  //                                    .txd
	);

	wire         altpll_clks_c0_clk;                                            // ALTPLL_CLKS:c0 -> [EXT_SDRAM_PROGMEM:clk, GPI0_BUTN:clk, GPI1_DIPSW:clk, GPO2_LEDG:clk, JTAG_UART_DBG:clk, NIOSV_M_CPU:clk, SOC_SYSID:clock, UART_SERIAL_COM:clk, irq_mapper:clk, irq_synchronizer:sender_clk, mm_interconnect_0:ALTPLL_CLKS_c0_clk, rst_controller_001:clk]
	wire         altpll_clks_c2_clk;                                            // ALTPLL_CLKS:c2 -> [EPCS_FLASH_CONTROLLER:clk, irq_synchronizer:receiver_clk, mm_interconnect_0:ALTPLL_CLKS_c2_clk, rst_controller:clk]
	wire  [31:0] niosv_m_cpu_data_manager_awaddr;                               // NIOSV_M_CPU:data_manager_awaddr -> mm_interconnect_0:NIOSV_M_CPU_data_manager_awaddr
	wire   [1:0] niosv_m_cpu_data_manager_bresp;                                // mm_interconnect_0:NIOSV_M_CPU_data_manager_bresp -> NIOSV_M_CPU:data_manager_bresp
	wire         niosv_m_cpu_data_manager_arready;                              // mm_interconnect_0:NIOSV_M_CPU_data_manager_arready -> NIOSV_M_CPU:data_manager_arready
	wire  [31:0] niosv_m_cpu_data_manager_rdata;                                // mm_interconnect_0:NIOSV_M_CPU_data_manager_rdata -> NIOSV_M_CPU:data_manager_rdata
	wire   [3:0] niosv_m_cpu_data_manager_wstrb;                                // NIOSV_M_CPU:data_manager_wstrb -> mm_interconnect_0:NIOSV_M_CPU_data_manager_wstrb
	wire         niosv_m_cpu_data_manager_wready;                               // mm_interconnect_0:NIOSV_M_CPU_data_manager_wready -> NIOSV_M_CPU:data_manager_wready
	wire         niosv_m_cpu_data_manager_awready;                              // mm_interconnect_0:NIOSV_M_CPU_data_manager_awready -> NIOSV_M_CPU:data_manager_awready
	wire         niosv_m_cpu_data_manager_rready;                               // NIOSV_M_CPU:data_manager_rready -> mm_interconnect_0:NIOSV_M_CPU_data_manager_rready
	wire         niosv_m_cpu_data_manager_bready;                               // NIOSV_M_CPU:data_manager_bready -> mm_interconnect_0:NIOSV_M_CPU_data_manager_bready
	wire         niosv_m_cpu_data_manager_wvalid;                               // NIOSV_M_CPU:data_manager_wvalid -> mm_interconnect_0:NIOSV_M_CPU_data_manager_wvalid
	wire  [31:0] niosv_m_cpu_data_manager_araddr;                               // NIOSV_M_CPU:data_manager_araddr -> mm_interconnect_0:NIOSV_M_CPU_data_manager_araddr
	wire   [2:0] niosv_m_cpu_data_manager_arprot;                               // NIOSV_M_CPU:data_manager_arprot -> mm_interconnect_0:NIOSV_M_CPU_data_manager_arprot
	wire   [1:0] niosv_m_cpu_data_manager_rresp;                                // mm_interconnect_0:NIOSV_M_CPU_data_manager_rresp -> NIOSV_M_CPU:data_manager_rresp
	wire   [2:0] niosv_m_cpu_data_manager_awprot;                               // NIOSV_M_CPU:data_manager_awprot -> mm_interconnect_0:NIOSV_M_CPU_data_manager_awprot
	wire  [31:0] niosv_m_cpu_data_manager_wdata;                                // NIOSV_M_CPU:data_manager_wdata -> mm_interconnect_0:NIOSV_M_CPU_data_manager_wdata
	wire         niosv_m_cpu_data_manager_arvalid;                              // NIOSV_M_CPU:data_manager_arvalid -> mm_interconnect_0:NIOSV_M_CPU_data_manager_arvalid
	wire         niosv_m_cpu_data_manager_bvalid;                               // mm_interconnect_0:NIOSV_M_CPU_data_manager_bvalid -> NIOSV_M_CPU:data_manager_bvalid
	wire         niosv_m_cpu_data_manager_awvalid;                              // NIOSV_M_CPU:data_manager_awvalid -> mm_interconnect_0:NIOSV_M_CPU_data_manager_awvalid
	wire         niosv_m_cpu_data_manager_rvalid;                               // mm_interconnect_0:NIOSV_M_CPU_data_manager_rvalid -> NIOSV_M_CPU:data_manager_rvalid
	wire  [31:0] niosv_m_cpu_instruction_manager_awaddr;                        // NIOSV_M_CPU:instruction_manager_awaddr -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_awaddr
	wire   [1:0] niosv_m_cpu_instruction_manager_bresp;                         // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_bresp -> NIOSV_M_CPU:instruction_manager_bresp
	wire         niosv_m_cpu_instruction_manager_arready;                       // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_arready -> NIOSV_M_CPU:instruction_manager_arready
	wire  [31:0] niosv_m_cpu_instruction_manager_rdata;                         // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_rdata -> NIOSV_M_CPU:instruction_manager_rdata
	wire   [3:0] niosv_m_cpu_instruction_manager_wstrb;                         // NIOSV_M_CPU:instruction_manager_wstrb -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_wstrb
	wire         niosv_m_cpu_instruction_manager_wready;                        // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_wready -> NIOSV_M_CPU:instruction_manager_wready
	wire         niosv_m_cpu_instruction_manager_awready;                       // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_awready -> NIOSV_M_CPU:instruction_manager_awready
	wire         niosv_m_cpu_instruction_manager_rready;                        // NIOSV_M_CPU:instruction_manager_rready -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_rready
	wire         niosv_m_cpu_instruction_manager_bready;                        // NIOSV_M_CPU:instruction_manager_bready -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_bready
	wire         niosv_m_cpu_instruction_manager_wvalid;                        // NIOSV_M_CPU:instruction_manager_wvalid -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_wvalid
	wire  [31:0] niosv_m_cpu_instruction_manager_araddr;                        // NIOSV_M_CPU:instruction_manager_araddr -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_araddr
	wire   [2:0] niosv_m_cpu_instruction_manager_arprot;                        // NIOSV_M_CPU:instruction_manager_arprot -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_arprot
	wire   [1:0] niosv_m_cpu_instruction_manager_rresp;                         // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_rresp -> NIOSV_M_CPU:instruction_manager_rresp
	wire   [2:0] niosv_m_cpu_instruction_manager_awprot;                        // NIOSV_M_CPU:instruction_manager_awprot -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_awprot
	wire  [31:0] niosv_m_cpu_instruction_manager_wdata;                         // NIOSV_M_CPU:instruction_manager_wdata -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_wdata
	wire         niosv_m_cpu_instruction_manager_arvalid;                       // NIOSV_M_CPU:instruction_manager_arvalid -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_arvalid
	wire         niosv_m_cpu_instruction_manager_bvalid;                        // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_bvalid -> NIOSV_M_CPU:instruction_manager_bvalid
	wire         niosv_m_cpu_instruction_manager_awvalid;                       // NIOSV_M_CPU:instruction_manager_awvalid -> mm_interconnect_0:NIOSV_M_CPU_instruction_manager_awvalid
	wire         niosv_m_cpu_instruction_manager_rvalid;                        // mm_interconnect_0:NIOSV_M_CPU_instruction_manager_rvalid -> NIOSV_M_CPU:instruction_manager_rvalid
	wire         mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_chipselect -> JTAG_UART_DBG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_readdata;    // JTAG_UART_DBG:av_readdata -> mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_waitrequest; // JTAG_UART_DBG:av_waitrequest -> mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_address -> JTAG_UART_DBG:av_address
	wire         mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_read -> JTAG_UART_DBG:av_read_n
	wire         mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_write -> JTAG_UART_DBG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_UART_DBG_avalon_jtag_slave_writedata -> JTAG_UART_DBG:av_writedata
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_avl_csr_readdata;      // EPCS_FLASH_CONTROLLER:avl_csr_rddata -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_csr_readdata
	wire         mm_interconnect_0_epcs_flash_controller_avl_csr_waitrequest;   // EPCS_FLASH_CONTROLLER:avl_csr_waitrequest -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_csr_waitrequest
	wire   [2:0] mm_interconnect_0_epcs_flash_controller_avl_csr_address;       // mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_csr_address -> EPCS_FLASH_CONTROLLER:avl_csr_addr
	wire         mm_interconnect_0_epcs_flash_controller_avl_csr_read;          // mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_csr_read -> EPCS_FLASH_CONTROLLER:avl_csr_read
	wire         mm_interconnect_0_epcs_flash_controller_avl_csr_readdatavalid; // EPCS_FLASH_CONTROLLER:avl_csr_rddata_valid -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_csr_readdatavalid
	wire         mm_interconnect_0_epcs_flash_controller_avl_csr_write;         // mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_csr_write -> EPCS_FLASH_CONTROLLER:avl_csr_write
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_avl_csr_writedata;     // mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_csr_writedata -> EPCS_FLASH_CONTROLLER:avl_csr_wrdata
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_avl_mem_readdata;      // EPCS_FLASH_CONTROLLER:avl_mem_rddata -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_mem_readdata
	wire         mm_interconnect_0_epcs_flash_controller_avl_mem_waitrequest;   // EPCS_FLASH_CONTROLLER:avl_mem_waitrequest -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_mem_waitrequest
	wire  [20:0] mm_interconnect_0_epcs_flash_controller_avl_mem_address;       // mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_mem_address -> EPCS_FLASH_CONTROLLER:avl_mem_addr
	wire         mm_interconnect_0_epcs_flash_controller_avl_mem_read;          // mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_mem_read -> EPCS_FLASH_CONTROLLER:avl_mem_read
	wire   [3:0] mm_interconnect_0_epcs_flash_controller_avl_mem_byteenable;    // mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_mem_byteenable -> EPCS_FLASH_CONTROLLER:avl_mem_byteenable
	wire         mm_interconnect_0_epcs_flash_controller_avl_mem_readdatavalid; // EPCS_FLASH_CONTROLLER:avl_mem_rddata_valid -> mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_mem_readdatavalid
	wire         mm_interconnect_0_epcs_flash_controller_avl_mem_write;         // mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_mem_write -> EPCS_FLASH_CONTROLLER:avl_mem_write
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_avl_mem_writedata;     // mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_mem_writedata -> EPCS_FLASH_CONTROLLER:avl_mem_wrdata
	wire   [6:0] mm_interconnect_0_epcs_flash_controller_avl_mem_burstcount;    // mm_interconnect_0:EPCS_FLASH_CONTROLLER_avl_mem_burstcount -> EPCS_FLASH_CONTROLLER:avl_mem_burstcount
	wire  [31:0] mm_interconnect_0_soc_sysid_control_slave_readdata;            // SOC_SYSID:readdata -> mm_interconnect_0:SOC_SYSID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_soc_sysid_control_slave_address;             // mm_interconnect_0:SOC_SYSID_control_slave_address -> SOC_SYSID:address
	wire  [31:0] mm_interconnect_0_niosv_m_cpu_dm_agent_readdata;               // NIOSV_M_CPU:dm_agent_readdata -> mm_interconnect_0:NIOSV_M_CPU_dm_agent_readdata
	wire         mm_interconnect_0_niosv_m_cpu_dm_agent_waitrequest;            // NIOSV_M_CPU:dm_agent_waitrequest -> mm_interconnect_0:NIOSV_M_CPU_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_niosv_m_cpu_dm_agent_address;                // mm_interconnect_0:NIOSV_M_CPU_dm_agent_address -> NIOSV_M_CPU:dm_agent_address
	wire         mm_interconnect_0_niosv_m_cpu_dm_agent_read;                   // mm_interconnect_0:NIOSV_M_CPU_dm_agent_read -> NIOSV_M_CPU:dm_agent_read
	wire         mm_interconnect_0_niosv_m_cpu_dm_agent_readdatavalid;          // NIOSV_M_CPU:dm_agent_readdatavalid -> mm_interconnect_0:NIOSV_M_CPU_dm_agent_readdatavalid
	wire         mm_interconnect_0_niosv_m_cpu_dm_agent_write;                  // mm_interconnect_0:NIOSV_M_CPU_dm_agent_write -> NIOSV_M_CPU:dm_agent_write
	wire  [31:0] mm_interconnect_0_niosv_m_cpu_dm_agent_writedata;              // mm_interconnect_0:NIOSV_M_CPU_dm_agent_writedata -> NIOSV_M_CPU:dm_agent_writedata
	wire  [31:0] mm_interconnect_0_altpll_clks_pll_slave_readdata;              // ALTPLL_CLKS:readdata -> mm_interconnect_0:ALTPLL_CLKS_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_clks_pll_slave_address;               // mm_interconnect_0:ALTPLL_CLKS_pll_slave_address -> ALTPLL_CLKS:address
	wire         mm_interconnect_0_altpll_clks_pll_slave_read;                  // mm_interconnect_0:ALTPLL_CLKS_pll_slave_read -> ALTPLL_CLKS:read
	wire         mm_interconnect_0_altpll_clks_pll_slave_write;                 // mm_interconnect_0:ALTPLL_CLKS_pll_slave_write -> ALTPLL_CLKS:write
	wire  [31:0] mm_interconnect_0_altpll_clks_pll_slave_writedata;             // mm_interconnect_0:ALTPLL_CLKS_pll_slave_writedata -> ALTPLL_CLKS:writedata
	wire         mm_interconnect_0_uart_serial_com_s1_chipselect;               // mm_interconnect_0:UART_SERIAL_COM_s1_chipselect -> UART_SERIAL_COM:chipselect
	wire  [15:0] mm_interconnect_0_uart_serial_com_s1_readdata;                 // UART_SERIAL_COM:readdata -> mm_interconnect_0:UART_SERIAL_COM_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_serial_com_s1_address;                  // mm_interconnect_0:UART_SERIAL_COM_s1_address -> UART_SERIAL_COM:address
	wire         mm_interconnect_0_uart_serial_com_s1_read;                     // mm_interconnect_0:UART_SERIAL_COM_s1_read -> UART_SERIAL_COM:read_n
	wire         mm_interconnect_0_uart_serial_com_s1_begintransfer;            // mm_interconnect_0:UART_SERIAL_COM_s1_begintransfer -> UART_SERIAL_COM:begintransfer
	wire         mm_interconnect_0_uart_serial_com_s1_write;                    // mm_interconnect_0:UART_SERIAL_COM_s1_write -> UART_SERIAL_COM:write_n
	wire  [15:0] mm_interconnect_0_uart_serial_com_s1_writedata;                // mm_interconnect_0:UART_SERIAL_COM_s1_writedata -> UART_SERIAL_COM:writedata
	wire         mm_interconnect_0_gpi0_butn_s1_chipselect;                     // mm_interconnect_0:GPI0_BUTN_s1_chipselect -> GPI0_BUTN:chipselect
	wire  [31:0] mm_interconnect_0_gpi0_butn_s1_readdata;                       // GPI0_BUTN:readdata -> mm_interconnect_0:GPI0_BUTN_s1_readdata
	wire   [1:0] mm_interconnect_0_gpi0_butn_s1_address;                        // mm_interconnect_0:GPI0_BUTN_s1_address -> GPI0_BUTN:address
	wire         mm_interconnect_0_gpi0_butn_s1_write;                          // mm_interconnect_0:GPI0_BUTN_s1_write -> GPI0_BUTN:write_n
	wire  [31:0] mm_interconnect_0_gpi0_butn_s1_writedata;                      // mm_interconnect_0:GPI0_BUTN_s1_writedata -> GPI0_BUTN:writedata
	wire         mm_interconnect_0_gpi1_dipsw_s1_chipselect;                    // mm_interconnect_0:GPI1_DIPSW_s1_chipselect -> GPI1_DIPSW:chipselect
	wire  [31:0] mm_interconnect_0_gpi1_dipsw_s1_readdata;                      // GPI1_DIPSW:readdata -> mm_interconnect_0:GPI1_DIPSW_s1_readdata
	wire   [1:0] mm_interconnect_0_gpi1_dipsw_s1_address;                       // mm_interconnect_0:GPI1_DIPSW_s1_address -> GPI1_DIPSW:address
	wire         mm_interconnect_0_gpi1_dipsw_s1_write;                         // mm_interconnect_0:GPI1_DIPSW_s1_write -> GPI1_DIPSW:write_n
	wire  [31:0] mm_interconnect_0_gpi1_dipsw_s1_writedata;                     // mm_interconnect_0:GPI1_DIPSW_s1_writedata -> GPI1_DIPSW:writedata
	wire         mm_interconnect_0_gpo2_ledg_s1_chipselect;                     // mm_interconnect_0:GPO2_LEDG_s1_chipselect -> GPO2_LEDG:chipselect
	wire  [31:0] mm_interconnect_0_gpo2_ledg_s1_readdata;                       // GPO2_LEDG:readdata -> mm_interconnect_0:GPO2_LEDG_s1_readdata
	wire   [2:0] mm_interconnect_0_gpo2_ledg_s1_address;                        // mm_interconnect_0:GPO2_LEDG_s1_address -> GPO2_LEDG:address
	wire         mm_interconnect_0_gpo2_ledg_s1_write;                          // mm_interconnect_0:GPO2_LEDG_s1_write -> GPO2_LEDG:write_n
	wire  [31:0] mm_interconnect_0_gpo2_ledg_s1_writedata;                      // mm_interconnect_0:GPO2_LEDG_s1_writedata -> GPO2_LEDG:writedata
	wire         mm_interconnect_0_ext_sdram_progmem_s1_chipselect;             // mm_interconnect_0:EXT_SDRAM_PROGMEM_s1_chipselect -> EXT_SDRAM_PROGMEM:az_cs
	wire  [15:0] mm_interconnect_0_ext_sdram_progmem_s1_readdata;               // EXT_SDRAM_PROGMEM:za_data -> mm_interconnect_0:EXT_SDRAM_PROGMEM_s1_readdata
	wire         mm_interconnect_0_ext_sdram_progmem_s1_waitrequest;            // EXT_SDRAM_PROGMEM:za_waitrequest -> mm_interconnect_0:EXT_SDRAM_PROGMEM_s1_waitrequest
	wire  [23:0] mm_interconnect_0_ext_sdram_progmem_s1_address;                // mm_interconnect_0:EXT_SDRAM_PROGMEM_s1_address -> EXT_SDRAM_PROGMEM:az_addr
	wire         mm_interconnect_0_ext_sdram_progmem_s1_read;                   // mm_interconnect_0:EXT_SDRAM_PROGMEM_s1_read -> EXT_SDRAM_PROGMEM:az_rd_n
	wire   [1:0] mm_interconnect_0_ext_sdram_progmem_s1_byteenable;             // mm_interconnect_0:EXT_SDRAM_PROGMEM_s1_byteenable -> EXT_SDRAM_PROGMEM:az_be_n
	wire         mm_interconnect_0_ext_sdram_progmem_s1_readdatavalid;          // EXT_SDRAM_PROGMEM:za_valid -> mm_interconnect_0:EXT_SDRAM_PROGMEM_s1_readdatavalid
	wire         mm_interconnect_0_ext_sdram_progmem_s1_write;                  // mm_interconnect_0:EXT_SDRAM_PROGMEM_s1_write -> EXT_SDRAM_PROGMEM:az_wr_n
	wire  [15:0] mm_interconnect_0_ext_sdram_progmem_s1_writedata;              // mm_interconnect_0:EXT_SDRAM_PROGMEM_s1_writedata -> EXT_SDRAM_PROGMEM:az_data
	wire  [31:0] mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdata;         // NIOSV_M_CPU:timer_sw_agent_readdata -> mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_readdata
	wire         mm_interconnect_0_niosv_m_cpu_timer_sw_agent_waitrequest;      // NIOSV_M_CPU:timer_sw_agent_waitrequest -> mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_waitrequest
	wire   [5:0] mm_interconnect_0_niosv_m_cpu_timer_sw_agent_address;          // mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_address -> NIOSV_M_CPU:timer_sw_agent_address
	wire         mm_interconnect_0_niosv_m_cpu_timer_sw_agent_read;             // mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_read -> NIOSV_M_CPU:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_niosv_m_cpu_timer_sw_agent_byteenable;       // mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_byteenable -> NIOSV_M_CPU:timer_sw_agent_byteenable
	wire         mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdatavalid;    // NIOSV_M_CPU:timer_sw_agent_readdatavalid -> mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_niosv_m_cpu_timer_sw_agent_write;            // mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_write -> NIOSV_M_CPU:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_niosv_m_cpu_timer_sw_agent_writedata;        // mm_interconnect_0:NIOSV_M_CPU_timer_sw_agent_writedata -> NIOSV_M_CPU:timer_sw_agent_writedata
	wire         irq_mapper_receiver1_irq;                                      // JTAG_UART_DBG:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                      // UART_SERIAL_COM:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                      // GPI0_BUTN:irq -> irq_mapper:receiver3_irq
	wire  [15:0] niosv_m_cpu_platform_irq_rx_irq;                               // irq_mapper:sender_irq -> NIOSV_M_CPU:platform_irq_rx_irq
	wire         irq_mapper_receiver0_irq;                                      // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                 // EPCS_FLASH_CONTROLLER:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [EPCS_FLASH_CONTROLLER:reset_n, irq_synchronizer:receiver_reset, mm_interconnect_0:EPCS_FLASH_CONTROLLER_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [EXT_SDRAM_PROGMEM:reset_n, GPI0_BUTN:reset_n, GPI1_DIPSW:reset_n, GPO2_LEDG:reset_n, JTAG_UART_DBG:rst_n, NIOSV_M_CPU:reset_reset, SOC_SYSID:reset_n, UART_SERIAL_COM:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:NIOSV_M_CPU_reset_reset_bridge_in_reset_reset]

	NIOSV_SOC_ALTPLL_CLKS altpll_clks (
		.clk                (in_clock_bridge_clk_clk),                           //       inclk_interface.clk
		.reset              (~in_reset_bridge_reset_reset_n),                    // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_clks_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_clks_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_clks_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_clks_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_clks_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_clks_c0_clk),                                //                    c0.clk
		.c1                 (altpll_clks_sdram_clk_clk),                         //                    c1.clk
		.c2                 (altpll_clks_c2_clk),                                //                    c2.clk
		.areset             (altpll_clks_areset_in_export),                      //        areset_conduit.export
		.locked             (altpll_clks_locked_out_export),                     //        locked_conduit.export
		.scandone           (),                                                  //           (terminated)
		.scandataout        (),                                                  //           (terminated)
		.phasedone          (),                                                  //           (terminated)
		.phasecounterselect (4'b0000),                                           //           (terminated)
		.phaseupdown        (1'b0),                                              //           (terminated)
		.phasestep          (1'b0),                                              //           (terminated)
		.scanclk            (1'b0),                                              //           (terminated)
		.scanclkena         (1'b0),                                              //           (terminated)
		.scandata           (1'b0),                                              //           (terminated)
		.configupdate       (1'b0)                                               //           (terminated)
	);

	NIOSV_SOC_EPCS_FLASH_CONTROLLER #(
		.DEVICE_FAMILY     ("Cyclone IV E"),
		.ASI_WIDTH         (1),
		.CS_WIDTH          (1),
		.ADDR_WIDTH        (21),
		.ASMI_ADDR_WIDTH   (24),
		.ENABLE_4BYTE_ADDR (0),
		.CHIP_SELS         (1)
	) epcs_flash_controller (
		.clk                  (altpll_clks_c2_clk),                                            //       clock_sink.clk
		.reset_n              (~rst_controller_reset_out_reset),                               //            reset.reset_n
		.avl_csr_read         (mm_interconnect_0_epcs_flash_controller_avl_csr_read),          //          avl_csr.read
		.avl_csr_waitrequest  (mm_interconnect_0_epcs_flash_controller_avl_csr_waitrequest),   //                 .waitrequest
		.avl_csr_write        (mm_interconnect_0_epcs_flash_controller_avl_csr_write),         //                 .write
		.avl_csr_addr         (mm_interconnect_0_epcs_flash_controller_avl_csr_address),       //                 .address
		.avl_csr_wrdata       (mm_interconnect_0_epcs_flash_controller_avl_csr_writedata),     //                 .writedata
		.avl_csr_rddata       (mm_interconnect_0_epcs_flash_controller_avl_csr_readdata),      //                 .readdata
		.avl_csr_rddata_valid (mm_interconnect_0_epcs_flash_controller_avl_csr_readdatavalid), //                 .readdatavalid
		.avl_mem_write        (mm_interconnect_0_epcs_flash_controller_avl_mem_write),         //          avl_mem.write
		.avl_mem_burstcount   (mm_interconnect_0_epcs_flash_controller_avl_mem_burstcount),    //                 .burstcount
		.avl_mem_waitrequest  (mm_interconnect_0_epcs_flash_controller_avl_mem_waitrequest),   //                 .waitrequest
		.avl_mem_read         (mm_interconnect_0_epcs_flash_controller_avl_mem_read),          //                 .read
		.avl_mem_addr         (mm_interconnect_0_epcs_flash_controller_avl_mem_address),       //                 .address
		.avl_mem_wrdata       (mm_interconnect_0_epcs_flash_controller_avl_mem_writedata),     //                 .writedata
		.avl_mem_rddata       (mm_interconnect_0_epcs_flash_controller_avl_mem_readdata),      //                 .readdata
		.avl_mem_rddata_valid (mm_interconnect_0_epcs_flash_controller_avl_mem_readdatavalid), //                 .readdatavalid
		.avl_mem_byteenable   (mm_interconnect_0_epcs_flash_controller_avl_mem_byteenable),    //                 .byteenable
		.irq                  (irq_synchronizer_receiver_irq)                                  // interrupt_sender.irq
	);

	NIOSV_SOC_EXT_SDRAM_PROGMEM ext_sdram_progmem (
		.clk            (altpll_clks_c0_clk),                                   //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                  // reset.reset_n
		.az_addr        (mm_interconnect_0_ext_sdram_progmem_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_ext_sdram_progmem_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_ext_sdram_progmem_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_ext_sdram_progmem_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_ext_sdram_progmem_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_ext_sdram_progmem_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_ext_sdram_progmem_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_ext_sdram_progmem_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_ext_sdram_progmem_s1_waitrequest),   //      .waitrequest
		.zs_addr        (ext_sdram_progmem_wire_addr),                          //  wire.export
		.zs_ba          (ext_sdram_progmem_wire_ba),                            //      .export
		.zs_cas_n       (ext_sdram_progmem_wire_cas_n),                         //      .export
		.zs_cke         (ext_sdram_progmem_wire_cke),                           //      .export
		.zs_cs_n        (ext_sdram_progmem_wire_cs_n),                          //      .export
		.zs_dq          (ext_sdram_progmem_wire_dq),                            //      .export
		.zs_dqm         (ext_sdram_progmem_wire_dqm),                           //      .export
		.zs_ras_n       (ext_sdram_progmem_wire_ras_n),                         //      .export
		.zs_we_n        (ext_sdram_progmem_wire_we_n)                           //      .export
	);

	NIOSV_SOC_GPI0_BUTN gpi0_butn (
		.clk        (altpll_clks_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_gpi0_butn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpi0_butn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpi0_butn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpi0_butn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpi0_butn_s1_readdata),   //                    .readdata
		.in_port    (gpi0_butn_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                   //                 irq.irq
	);

	NIOSV_SOC_GPI1_DIPSW gpi1_dipsw (
		.clk        (altpll_clks_c0_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_gpi1_dipsw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpi1_dipsw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpi1_dipsw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpi1_dipsw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpi1_dipsw_s1_readdata),   //                    .readdata
		.in_port    (gpi1_dipsw_external_connection_export)       // external_connection.export
	);

	NIOSV_SOC_GPO2_LEDG gpo2_ledg (
		.clk        (altpll_clks_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_gpo2_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpo2_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpo2_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpo2_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpo2_ledg_s1_readdata),   //                    .readdata
		.out_port   (gpo2_ledg_external_connection_export)       // external_connection.export
	);

	NIOSV_SOC_JTAG_UART_DBG jtag_uart_dbg (
		.clk            (altpll_clks_c0_clk),                                            //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                       //               irq.irq
	);

	NIOSV_SOC_NIOSV_M_CPU niosv_m_cpu (
		.clk                          (altpll_clks_c0_clk),                                         //                 clk.clk
		.reset_reset                  (rst_controller_001_reset_out_reset),                         //               reset.reset
		.platform_irq_rx_irq          (niosv_m_cpu_platform_irq_rx_irq),                            //     platform_irq_rx.irq
		.timer_sw_agent_write         (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_write),         //      timer_sw_agent.write
		.timer_sw_agent_writedata     (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_writedata),     //                    .writedata
		.timer_sw_agent_byteenable    (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_byteenable),    //                    .byteenable
		.timer_sw_agent_address       (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_address),       //                    .address
		.timer_sw_agent_read          (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_read),          //                    .read
		.timer_sw_agent_readdata      (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdata),      //                    .readdata
		.timer_sw_agent_readdatavalid (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdatavalid), //                    .readdatavalid
		.timer_sw_agent_waitrequest   (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_waitrequest),   //                    .waitrequest
		.instruction_manager_awaddr   (niosv_m_cpu_instruction_manager_awaddr),                     // instruction_manager.awaddr
		.instruction_manager_awprot   (niosv_m_cpu_instruction_manager_awprot),                     //                    .awprot
		.instruction_manager_awvalid  (niosv_m_cpu_instruction_manager_awvalid),                    //                    .awvalid
		.instruction_manager_awready  (niosv_m_cpu_instruction_manager_awready),                    //                    .awready
		.instruction_manager_wdata    (niosv_m_cpu_instruction_manager_wdata),                      //                    .wdata
		.instruction_manager_wstrb    (niosv_m_cpu_instruction_manager_wstrb),                      //                    .wstrb
		.instruction_manager_wvalid   (niosv_m_cpu_instruction_manager_wvalid),                     //                    .wvalid
		.instruction_manager_wready   (niosv_m_cpu_instruction_manager_wready),                     //                    .wready
		.instruction_manager_bresp    (niosv_m_cpu_instruction_manager_bresp),                      //                    .bresp
		.instruction_manager_bvalid   (niosv_m_cpu_instruction_manager_bvalid),                     //                    .bvalid
		.instruction_manager_bready   (niosv_m_cpu_instruction_manager_bready),                     //                    .bready
		.instruction_manager_araddr   (niosv_m_cpu_instruction_manager_araddr),                     //                    .araddr
		.instruction_manager_arprot   (niosv_m_cpu_instruction_manager_arprot),                     //                    .arprot
		.instruction_manager_arvalid  (niosv_m_cpu_instruction_manager_arvalid),                    //                    .arvalid
		.instruction_manager_arready  (niosv_m_cpu_instruction_manager_arready),                    //                    .arready
		.instruction_manager_rdata    (niosv_m_cpu_instruction_manager_rdata),                      //                    .rdata
		.instruction_manager_rresp    (niosv_m_cpu_instruction_manager_rresp),                      //                    .rresp
		.instruction_manager_rvalid   (niosv_m_cpu_instruction_manager_rvalid),                     //                    .rvalid
		.instruction_manager_rready   (niosv_m_cpu_instruction_manager_rready),                     //                    .rready
		.data_manager_awaddr          (niosv_m_cpu_data_manager_awaddr),                            //        data_manager.awaddr
		.data_manager_awprot          (niosv_m_cpu_data_manager_awprot),                            //                    .awprot
		.data_manager_awvalid         (niosv_m_cpu_data_manager_awvalid),                           //                    .awvalid
		.data_manager_awready         (niosv_m_cpu_data_manager_awready),                           //                    .awready
		.data_manager_wdata           (niosv_m_cpu_data_manager_wdata),                             //                    .wdata
		.data_manager_wstrb           (niosv_m_cpu_data_manager_wstrb),                             //                    .wstrb
		.data_manager_wvalid          (niosv_m_cpu_data_manager_wvalid),                            //                    .wvalid
		.data_manager_wready          (niosv_m_cpu_data_manager_wready),                            //                    .wready
		.data_manager_bresp           (niosv_m_cpu_data_manager_bresp),                             //                    .bresp
		.data_manager_bvalid          (niosv_m_cpu_data_manager_bvalid),                            //                    .bvalid
		.data_manager_bready          (niosv_m_cpu_data_manager_bready),                            //                    .bready
		.data_manager_araddr          (niosv_m_cpu_data_manager_araddr),                            //                    .araddr
		.data_manager_arprot          (niosv_m_cpu_data_manager_arprot),                            //                    .arprot
		.data_manager_arvalid         (niosv_m_cpu_data_manager_arvalid),                           //                    .arvalid
		.data_manager_arready         (niosv_m_cpu_data_manager_arready),                           //                    .arready
		.data_manager_rdata           (niosv_m_cpu_data_manager_rdata),                             //                    .rdata
		.data_manager_rresp           (niosv_m_cpu_data_manager_rresp),                             //                    .rresp
		.data_manager_rvalid          (niosv_m_cpu_data_manager_rvalid),                            //                    .rvalid
		.data_manager_rready          (niosv_m_cpu_data_manager_rready),                            //                    .rready
		.dm_agent_write               (mm_interconnect_0_niosv_m_cpu_dm_agent_write),               //            dm_agent.write
		.dm_agent_writedata           (mm_interconnect_0_niosv_m_cpu_dm_agent_writedata),           //                    .writedata
		.dm_agent_address             (mm_interconnect_0_niosv_m_cpu_dm_agent_address),             //                    .address
		.dm_agent_read                (mm_interconnect_0_niosv_m_cpu_dm_agent_read),                //                    .read
		.dm_agent_readdata            (mm_interconnect_0_niosv_m_cpu_dm_agent_readdata),            //                    .readdata
		.dm_agent_readdatavalid       (mm_interconnect_0_niosv_m_cpu_dm_agent_readdatavalid),       //                    .readdatavalid
		.dm_agent_waitrequest         (mm_interconnect_0_niosv_m_cpu_dm_agent_waitrequest),         //                    .waitrequest
		.cpu_ecc_status_ecc_status    (),                                                           //      cpu_ecc_status.ecc_status
		.cpu_ecc_status_ecc_source    ()                                                            //                    .ecc_source
	);

	NIOSV_SOC_SOC_SYSID soc_sysid (
		.clock    (altpll_clks_c0_clk),                                 //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_soc_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_soc_sysid_control_slave_address)   //              .address
	);

	NIOSV_SOC_UART_SERIAL_COM uart_serial_com (
		.clk           (altpll_clks_c0_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                //               reset.reset_n
		.address       (mm_interconnect_0_uart_serial_com_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_serial_com_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_serial_com_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_serial_com_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_serial_com_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_serial_com_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_serial_com_s1_readdata),      //                    .readdata
		.rxd           (uart_serial_com_external_connection_rxd),            // external_connection.export
		.txd           (uart_serial_com_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver2_irq)                            //                 irq.irq
	);

	NIOSV_SOC_mm_interconnect_0 mm_interconnect_0 (
		.NIOSV_M_CPU_data_manager_awaddr                               (niosv_m_cpu_data_manager_awaddr),                               //                                NIOSV_M_CPU_data_manager.awaddr
		.NIOSV_M_CPU_data_manager_awprot                               (niosv_m_cpu_data_manager_awprot),                               //                                                        .awprot
		.NIOSV_M_CPU_data_manager_awvalid                              (niosv_m_cpu_data_manager_awvalid),                              //                                                        .awvalid
		.NIOSV_M_CPU_data_manager_awready                              (niosv_m_cpu_data_manager_awready),                              //                                                        .awready
		.NIOSV_M_CPU_data_manager_wdata                                (niosv_m_cpu_data_manager_wdata),                                //                                                        .wdata
		.NIOSV_M_CPU_data_manager_wstrb                                (niosv_m_cpu_data_manager_wstrb),                                //                                                        .wstrb
		.NIOSV_M_CPU_data_manager_wvalid                               (niosv_m_cpu_data_manager_wvalid),                               //                                                        .wvalid
		.NIOSV_M_CPU_data_manager_wready                               (niosv_m_cpu_data_manager_wready),                               //                                                        .wready
		.NIOSV_M_CPU_data_manager_bresp                                (niosv_m_cpu_data_manager_bresp),                                //                                                        .bresp
		.NIOSV_M_CPU_data_manager_bvalid                               (niosv_m_cpu_data_manager_bvalid),                               //                                                        .bvalid
		.NIOSV_M_CPU_data_manager_bready                               (niosv_m_cpu_data_manager_bready),                               //                                                        .bready
		.NIOSV_M_CPU_data_manager_araddr                               (niosv_m_cpu_data_manager_araddr),                               //                                                        .araddr
		.NIOSV_M_CPU_data_manager_arprot                               (niosv_m_cpu_data_manager_arprot),                               //                                                        .arprot
		.NIOSV_M_CPU_data_manager_arvalid                              (niosv_m_cpu_data_manager_arvalid),                              //                                                        .arvalid
		.NIOSV_M_CPU_data_manager_arready                              (niosv_m_cpu_data_manager_arready),                              //                                                        .arready
		.NIOSV_M_CPU_data_manager_rdata                                (niosv_m_cpu_data_manager_rdata),                                //                                                        .rdata
		.NIOSV_M_CPU_data_manager_rresp                                (niosv_m_cpu_data_manager_rresp),                                //                                                        .rresp
		.NIOSV_M_CPU_data_manager_rvalid                               (niosv_m_cpu_data_manager_rvalid),                               //                                                        .rvalid
		.NIOSV_M_CPU_data_manager_rready                               (niosv_m_cpu_data_manager_rready),                               //                                                        .rready
		.NIOSV_M_CPU_instruction_manager_awaddr                        (niosv_m_cpu_instruction_manager_awaddr),                        //                         NIOSV_M_CPU_instruction_manager.awaddr
		.NIOSV_M_CPU_instruction_manager_awprot                        (niosv_m_cpu_instruction_manager_awprot),                        //                                                        .awprot
		.NIOSV_M_CPU_instruction_manager_awvalid                       (niosv_m_cpu_instruction_manager_awvalid),                       //                                                        .awvalid
		.NIOSV_M_CPU_instruction_manager_awready                       (niosv_m_cpu_instruction_manager_awready),                       //                                                        .awready
		.NIOSV_M_CPU_instruction_manager_wdata                         (niosv_m_cpu_instruction_manager_wdata),                         //                                                        .wdata
		.NIOSV_M_CPU_instruction_manager_wstrb                         (niosv_m_cpu_instruction_manager_wstrb),                         //                                                        .wstrb
		.NIOSV_M_CPU_instruction_manager_wvalid                        (niosv_m_cpu_instruction_manager_wvalid),                        //                                                        .wvalid
		.NIOSV_M_CPU_instruction_manager_wready                        (niosv_m_cpu_instruction_manager_wready),                        //                                                        .wready
		.NIOSV_M_CPU_instruction_manager_bresp                         (niosv_m_cpu_instruction_manager_bresp),                         //                                                        .bresp
		.NIOSV_M_CPU_instruction_manager_bvalid                        (niosv_m_cpu_instruction_manager_bvalid),                        //                                                        .bvalid
		.NIOSV_M_CPU_instruction_manager_bready                        (niosv_m_cpu_instruction_manager_bready),                        //                                                        .bready
		.NIOSV_M_CPU_instruction_manager_araddr                        (niosv_m_cpu_instruction_manager_araddr),                        //                                                        .araddr
		.NIOSV_M_CPU_instruction_manager_arprot                        (niosv_m_cpu_instruction_manager_arprot),                        //                                                        .arprot
		.NIOSV_M_CPU_instruction_manager_arvalid                       (niosv_m_cpu_instruction_manager_arvalid),                       //                                                        .arvalid
		.NIOSV_M_CPU_instruction_manager_arready                       (niosv_m_cpu_instruction_manager_arready),                       //                                                        .arready
		.NIOSV_M_CPU_instruction_manager_rdata                         (niosv_m_cpu_instruction_manager_rdata),                         //                                                        .rdata
		.NIOSV_M_CPU_instruction_manager_rresp                         (niosv_m_cpu_instruction_manager_rresp),                         //                                                        .rresp
		.NIOSV_M_CPU_instruction_manager_rvalid                        (niosv_m_cpu_instruction_manager_rvalid),                        //                                                        .rvalid
		.NIOSV_M_CPU_instruction_manager_rready                        (niosv_m_cpu_instruction_manager_rready),                        //                                                        .rready
		.ALTPLL_CLKS_c0_clk                                            (altpll_clks_c0_clk),                                            //                                          ALTPLL_CLKS_c0.clk
		.ALTPLL_CLKS_c2_clk                                            (altpll_clks_c2_clk),                                            //                                          ALTPLL_CLKS_c2.clk
		.IN_CLOCK_BRIDGE_out_clk_clk                                   (in_clock_bridge_clk_clk),                                       //                                 IN_CLOCK_BRIDGE_out_clk.clk
		.ALTPLL_CLKS_inclk_interface_reset_reset_bridge_in_reset_reset (~in_reset_bridge_reset_reset_n),                                // ALTPLL_CLKS_inclk_interface_reset_reset_bridge_in_reset.reset
		.EPCS_FLASH_CONTROLLER_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                                //       EPCS_FLASH_CONTROLLER_reset_reset_bridge_in_reset.reset
		.NIOSV_M_CPU_reset_reset_bridge_in_reset_reset                 (rst_controller_001_reset_out_reset),                            //                 NIOSV_M_CPU_reset_reset_bridge_in_reset.reset
		.ALTPLL_CLKS_pll_slave_address                                 (mm_interconnect_0_altpll_clks_pll_slave_address),               //                                   ALTPLL_CLKS_pll_slave.address
		.ALTPLL_CLKS_pll_slave_write                                   (mm_interconnect_0_altpll_clks_pll_slave_write),                 //                                                        .write
		.ALTPLL_CLKS_pll_slave_read                                    (mm_interconnect_0_altpll_clks_pll_slave_read),                  //                                                        .read
		.ALTPLL_CLKS_pll_slave_readdata                                (mm_interconnect_0_altpll_clks_pll_slave_readdata),              //                                                        .readdata
		.ALTPLL_CLKS_pll_slave_writedata                               (mm_interconnect_0_altpll_clks_pll_slave_writedata),             //                                                        .writedata
		.EPCS_FLASH_CONTROLLER_avl_csr_address                         (mm_interconnect_0_epcs_flash_controller_avl_csr_address),       //                           EPCS_FLASH_CONTROLLER_avl_csr.address
		.EPCS_FLASH_CONTROLLER_avl_csr_write                           (mm_interconnect_0_epcs_flash_controller_avl_csr_write),         //                                                        .write
		.EPCS_FLASH_CONTROLLER_avl_csr_read                            (mm_interconnect_0_epcs_flash_controller_avl_csr_read),          //                                                        .read
		.EPCS_FLASH_CONTROLLER_avl_csr_readdata                        (mm_interconnect_0_epcs_flash_controller_avl_csr_readdata),      //                                                        .readdata
		.EPCS_FLASH_CONTROLLER_avl_csr_writedata                       (mm_interconnect_0_epcs_flash_controller_avl_csr_writedata),     //                                                        .writedata
		.EPCS_FLASH_CONTROLLER_avl_csr_readdatavalid                   (mm_interconnect_0_epcs_flash_controller_avl_csr_readdatavalid), //                                                        .readdatavalid
		.EPCS_FLASH_CONTROLLER_avl_csr_waitrequest                     (mm_interconnect_0_epcs_flash_controller_avl_csr_waitrequest),   //                                                        .waitrequest
		.EPCS_FLASH_CONTROLLER_avl_mem_address                         (mm_interconnect_0_epcs_flash_controller_avl_mem_address),       //                           EPCS_FLASH_CONTROLLER_avl_mem.address
		.EPCS_FLASH_CONTROLLER_avl_mem_write                           (mm_interconnect_0_epcs_flash_controller_avl_mem_write),         //                                                        .write
		.EPCS_FLASH_CONTROLLER_avl_mem_read                            (mm_interconnect_0_epcs_flash_controller_avl_mem_read),          //                                                        .read
		.EPCS_FLASH_CONTROLLER_avl_mem_readdata                        (mm_interconnect_0_epcs_flash_controller_avl_mem_readdata),      //                                                        .readdata
		.EPCS_FLASH_CONTROLLER_avl_mem_writedata                       (mm_interconnect_0_epcs_flash_controller_avl_mem_writedata),     //                                                        .writedata
		.EPCS_FLASH_CONTROLLER_avl_mem_burstcount                      (mm_interconnect_0_epcs_flash_controller_avl_mem_burstcount),    //                                                        .burstcount
		.EPCS_FLASH_CONTROLLER_avl_mem_byteenable                      (mm_interconnect_0_epcs_flash_controller_avl_mem_byteenable),    //                                                        .byteenable
		.EPCS_FLASH_CONTROLLER_avl_mem_readdatavalid                   (mm_interconnect_0_epcs_flash_controller_avl_mem_readdatavalid), //                                                        .readdatavalid
		.EPCS_FLASH_CONTROLLER_avl_mem_waitrequest                     (mm_interconnect_0_epcs_flash_controller_avl_mem_waitrequest),   //                                                        .waitrequest
		.EXT_SDRAM_PROGMEM_s1_address                                  (mm_interconnect_0_ext_sdram_progmem_s1_address),                //                                    EXT_SDRAM_PROGMEM_s1.address
		.EXT_SDRAM_PROGMEM_s1_write                                    (mm_interconnect_0_ext_sdram_progmem_s1_write),                  //                                                        .write
		.EXT_SDRAM_PROGMEM_s1_read                                     (mm_interconnect_0_ext_sdram_progmem_s1_read),                   //                                                        .read
		.EXT_SDRAM_PROGMEM_s1_readdata                                 (mm_interconnect_0_ext_sdram_progmem_s1_readdata),               //                                                        .readdata
		.EXT_SDRAM_PROGMEM_s1_writedata                                (mm_interconnect_0_ext_sdram_progmem_s1_writedata),              //                                                        .writedata
		.EXT_SDRAM_PROGMEM_s1_byteenable                               (mm_interconnect_0_ext_sdram_progmem_s1_byteenable),             //                                                        .byteenable
		.EXT_SDRAM_PROGMEM_s1_readdatavalid                            (mm_interconnect_0_ext_sdram_progmem_s1_readdatavalid),          //                                                        .readdatavalid
		.EXT_SDRAM_PROGMEM_s1_waitrequest                              (mm_interconnect_0_ext_sdram_progmem_s1_waitrequest),            //                                                        .waitrequest
		.EXT_SDRAM_PROGMEM_s1_chipselect                               (mm_interconnect_0_ext_sdram_progmem_s1_chipselect),             //                                                        .chipselect
		.GPI0_BUTN_s1_address                                          (mm_interconnect_0_gpi0_butn_s1_address),                        //                                            GPI0_BUTN_s1.address
		.GPI0_BUTN_s1_write                                            (mm_interconnect_0_gpi0_butn_s1_write),                          //                                                        .write
		.GPI0_BUTN_s1_readdata                                         (mm_interconnect_0_gpi0_butn_s1_readdata),                       //                                                        .readdata
		.GPI0_BUTN_s1_writedata                                        (mm_interconnect_0_gpi0_butn_s1_writedata),                      //                                                        .writedata
		.GPI0_BUTN_s1_chipselect                                       (mm_interconnect_0_gpi0_butn_s1_chipselect),                     //                                                        .chipselect
		.GPI1_DIPSW_s1_address                                         (mm_interconnect_0_gpi1_dipsw_s1_address),                       //                                           GPI1_DIPSW_s1.address
		.GPI1_DIPSW_s1_write                                           (mm_interconnect_0_gpi1_dipsw_s1_write),                         //                                                        .write
		.GPI1_DIPSW_s1_readdata                                        (mm_interconnect_0_gpi1_dipsw_s1_readdata),                      //                                                        .readdata
		.GPI1_DIPSW_s1_writedata                                       (mm_interconnect_0_gpi1_dipsw_s1_writedata),                     //                                                        .writedata
		.GPI1_DIPSW_s1_chipselect                                      (mm_interconnect_0_gpi1_dipsw_s1_chipselect),                    //                                                        .chipselect
		.GPO2_LEDG_s1_address                                          (mm_interconnect_0_gpo2_ledg_s1_address),                        //                                            GPO2_LEDG_s1.address
		.GPO2_LEDG_s1_write                                            (mm_interconnect_0_gpo2_ledg_s1_write),                          //                                                        .write
		.GPO2_LEDG_s1_readdata                                         (mm_interconnect_0_gpo2_ledg_s1_readdata),                       //                                                        .readdata
		.GPO2_LEDG_s1_writedata                                        (mm_interconnect_0_gpo2_ledg_s1_writedata),                      //                                                        .writedata
		.GPO2_LEDG_s1_chipselect                                       (mm_interconnect_0_gpo2_ledg_s1_chipselect),                     //                                                        .chipselect
		.JTAG_UART_DBG_avalon_jtag_slave_address                       (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_address),     //                         JTAG_UART_DBG_avalon_jtag_slave.address
		.JTAG_UART_DBG_avalon_jtag_slave_write                         (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_write),       //                                                        .write
		.JTAG_UART_DBG_avalon_jtag_slave_read                          (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_read),        //                                                        .read
		.JTAG_UART_DBG_avalon_jtag_slave_readdata                      (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_readdata),    //                                                        .readdata
		.JTAG_UART_DBG_avalon_jtag_slave_writedata                     (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_writedata),   //                                                        .writedata
		.JTAG_UART_DBG_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_waitrequest), //                                                        .waitrequest
		.JTAG_UART_DBG_avalon_jtag_slave_chipselect                    (mm_interconnect_0_jtag_uart_dbg_avalon_jtag_slave_chipselect),  //                                                        .chipselect
		.NIOSV_M_CPU_dm_agent_address                                  (mm_interconnect_0_niosv_m_cpu_dm_agent_address),                //                                    NIOSV_M_CPU_dm_agent.address
		.NIOSV_M_CPU_dm_agent_write                                    (mm_interconnect_0_niosv_m_cpu_dm_agent_write),                  //                                                        .write
		.NIOSV_M_CPU_dm_agent_read                                     (mm_interconnect_0_niosv_m_cpu_dm_agent_read),                   //                                                        .read
		.NIOSV_M_CPU_dm_agent_readdata                                 (mm_interconnect_0_niosv_m_cpu_dm_agent_readdata),               //                                                        .readdata
		.NIOSV_M_CPU_dm_agent_writedata                                (mm_interconnect_0_niosv_m_cpu_dm_agent_writedata),              //                                                        .writedata
		.NIOSV_M_CPU_dm_agent_readdatavalid                            (mm_interconnect_0_niosv_m_cpu_dm_agent_readdatavalid),          //                                                        .readdatavalid
		.NIOSV_M_CPU_dm_agent_waitrequest                              (mm_interconnect_0_niosv_m_cpu_dm_agent_waitrequest),            //                                                        .waitrequest
		.NIOSV_M_CPU_timer_sw_agent_address                            (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_address),          //                              NIOSV_M_CPU_timer_sw_agent.address
		.NIOSV_M_CPU_timer_sw_agent_write                              (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_write),            //                                                        .write
		.NIOSV_M_CPU_timer_sw_agent_read                               (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_read),             //                                                        .read
		.NIOSV_M_CPU_timer_sw_agent_readdata                           (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdata),         //                                                        .readdata
		.NIOSV_M_CPU_timer_sw_agent_writedata                          (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_writedata),        //                                                        .writedata
		.NIOSV_M_CPU_timer_sw_agent_byteenable                         (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_byteenable),       //                                                        .byteenable
		.NIOSV_M_CPU_timer_sw_agent_readdatavalid                      (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_readdatavalid),    //                                                        .readdatavalid
		.NIOSV_M_CPU_timer_sw_agent_waitrequest                        (mm_interconnect_0_niosv_m_cpu_timer_sw_agent_waitrequest),      //                                                        .waitrequest
		.SOC_SYSID_control_slave_address                               (mm_interconnect_0_soc_sysid_control_slave_address),             //                                 SOC_SYSID_control_slave.address
		.SOC_SYSID_control_slave_readdata                              (mm_interconnect_0_soc_sysid_control_slave_readdata),            //                                                        .readdata
		.UART_SERIAL_COM_s1_address                                    (mm_interconnect_0_uart_serial_com_s1_address),                  //                                      UART_SERIAL_COM_s1.address
		.UART_SERIAL_COM_s1_write                                      (mm_interconnect_0_uart_serial_com_s1_write),                    //                                                        .write
		.UART_SERIAL_COM_s1_read                                       (mm_interconnect_0_uart_serial_com_s1_read),                     //                                                        .read
		.UART_SERIAL_COM_s1_readdata                                   (mm_interconnect_0_uart_serial_com_s1_readdata),                 //                                                        .readdata
		.UART_SERIAL_COM_s1_writedata                                  (mm_interconnect_0_uart_serial_com_s1_writedata),                //                                                        .writedata
		.UART_SERIAL_COM_s1_begintransfer                              (mm_interconnect_0_uart_serial_com_s1_begintransfer),            //                                                        .begintransfer
		.UART_SERIAL_COM_s1_chipselect                                 (mm_interconnect_0_uart_serial_com_s1_chipselect)                //                                                        .chipselect
	);

	NIOSV_SOC_irq_mapper irq_mapper (
		.clk           (altpll_clks_c0_clk),                 //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (niosv_m_cpu_platform_irq_rx_irq)     //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_clks_c2_clk),                 //       receiver_clk.clk
		.sender_clk     (altpll_clks_c0_clk),                 //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~in_reset_bridge_reset_reset_n), // reset_in0.reset
		.clk            (altpll_clks_c2_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~in_reset_bridge_reset_reset_n),     // reset_in0.reset
		.clk            (altpll_clks_c0_clk),                 //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
