��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��=�P��q�n'���}6𞆤m��j�I�� ۊ�E0��`� Sگ�v���ҢWs��[3 �z�XW��И n���W��PDo��Fس.<"t�bhS��A�P��M�5�I��mw?�h�s^,�O{ڕ�Ln��oA��!K9�2'�'�!W����̩Oٰ8��)��Ɉ|h�`O���se��
<C��x��o��c�`�'1�o#��+��	B
0�2O�I�2U�֛�n��ȵ��@�Ҭ�k�Yq�JVc�E&F�@��G�8�8�I�ܗO�[p��/�>���ţ�~}��J���u��^;X��R�UT��`�B��e֩�,�w� Mմ�'�F�P�8�5��T�Ԟ�C�đ��H%߂;h
,��'�A��%�8��_��� ���S
֚�� �V5�UÅZB�<�i�{ ~��-��M� s�hPO��k���"�۸9�ʉ�G���D�4��iXQ�"|r�8V��p�}J�"-�]��F/�(�)�Q���>��.,>[�]�|�b�E��sy��%�j���o;L#�t��`�?+֭�ySzT�^�,�]�HR�mZ���W��'���Z`�Ɓe�Jŗ�
X�c�'�R�u�!J�tW6{*5A�)E6�'S���u��t���/�?����o��}����i�n`\ƥ2Z
ݼI1O "���U�{v�fs��~������|B׫ۏ���$�r��d�f!�L؁�3�@3@4���E���������!�T�U�Ra��|y
�܌"3�"�����A-��M���c ��}?��(N0U.��2/�N�bz�I���I~�̀!yDP��r���[߸+���R���oߝS�F��J8�9sCP��T'�7�&��?G�uG8�{x������G�y�̸�Ur�+퉂d�~B{���-�l�1�܇���s�axcyMGl�!�S����\���us$�KIlv�^�>�j<$�a}v��[��F_��xR��$��_Dg�}���ǧ�]�l vE����2mD�h�7
�˦�0톝ZL��ʖ]tUD�"d�ft��}�_+#�Jc�#Q���׼%�{���C�ӼK�{T>A��]-#������)i\N
&.�@��7�1Ҋ�[t�T����G}�%i�*��J$z�U�}��J�tv�[nؔ��;��i�`��C�gP���Y�e�]���⨙���C?���*��1�:�M�8� z-�v yo�'fo�E�q�i�)�~�h�z|ma����Ѣ�q�Ֆ������H��V	&M;j���i���.]�~N�d�OȽ��f�wɾ�y�M�U+
*�
�mt��*��>
1ü�ja�^g��>��f�{SU��w���� M���{a_P.N��O����G�����QE���+N%A֐f�����ts�rS�&�Į<H/C�d	��b����o} J�O|�-����#������qx�q�Z��a��8{;ehc��(3�=v
*dK �ŷ�9��j2V�6��q��*PiFΗ�>3��p�8� ]�{N�W�[��|���@���K�ه�oo�����S1�Ę-�l]�����e
�|�R��`,�z�=���������.�ō�9�,kCA���q���J:e�b ��wF�q6�S"��>���1�l�U9���|�C+�9�^��:Qڞ��������结T��F*sN��n���7�t�ޗV�?u��:��3ӜC�b��\�d�&,r7�x��Z��;�[��=cx���&�9�W�ۂ(l���u�>��f�PX��82/�0J1ϵ�8���B��#f�-v/�kW��Č�-�sؾ�!)Z�C�X��0�iH{@���[�{�`ԥm����U��9(+k@�0b�P�S���˗� r̓�n���?�[��~.��٢hh�}f�k�vy�s��c%����+�4�O��<���]��x:���o)��$5\�`�i!��#��B	����N����/ַs�[{岨]���Y�RT��gU�������7�P׋J�[>O~?	9>|>?7 ]�ֵnD����%)ΔO���ą�`Sq�L���pZ�e��ɡ/�qV��hc��E�.w/8��!�^��W���?H��NH����S�t*����A�x����X�E|�j�A�sz��Vp%��y׮��������=���9�_�%��G�2� �,MPGJ\������Jd��E\�����NT�\{c�9da��D\l0���'&w�b?k
�m���v��/���C*�Hs�)�]P����Qg�y_<3!�NI#�����,���7���zP��4d5�'H1��!C��h�r��:�Q������^;���&٘�f��`�P
k��cF0|_]��p\��h��J۬w�w��5�	H��D+�8��BM��C�l����-��a7)�|�4a��k�Q��4���R��	J�;���{Q_��xF�����zԌ�#��6��}��aT�>��fyņըٱ^XT'������td�!5���*�	2�E���ơL�"��h�ٳ�^�@1��<�v�	*�2;�='���M2"�Q�q���\�L�ԭeY�;�v���#9���+c�M	yF�:�d���q����j#t�sLU��]�a_���2r4�)��F| je��F�#�O�MV�"1As#��K��w���xr���7ￓ��q>u$�gL�bK�f~<V�=?�4h�b�`+(��OSP�t�� ��t�j�f����i���a]�i�@�ْKV:m1!]�0	��=���X��!չl�/��y���ƛi6³}�yE�$/�mrۓ���xw�L7�8�3��hځ]�,��8!�PZ$h���
��y��S��z��e҆Y��F���>�E�ફp��s����V�E��߁tK?���3�yka�(�x�*Q�����������87�p�}��|g�N�#+�����vŏ�������2pb�ۆ-Tr�*��Mv�r�o�&6�J�F<QϬ��*2[\�k�͊l��L�"8H�����h�|��Nu	a�H� ^�5%%�o���/���ER!_�x��Ή�-m�mu$'ȷn��Bs+t�)zvU����P��8�t�|�҂�%AD��^�V4��6�}Ldz%����ɊO<�¥k4y�P1"�AE�\l|l�q�w�Mm��sݱz;�"*�9�n L&bY��S�C�qJ����ܩ�R�! 6�yj+w�_ $"��za��m�)$��ݾ��?]ݞC�Y6!�
m�D��㶍�8qq����ʍ�l�p��b��ٱ�����)$[N>z���J����YY�����<�I�	���s/�ꓰ�˂g�3� 4'�єA3T:Ϧlǥ�2}��\OS�	P�	�({m#�z{�ɯ#]CM��P>,�
��ȭ���,b� �����j9��[9F��p`a�'��7�}��T���A$��R���&,�w�LS.N�f�t$~���W�ks��w�X��̢ՔB���l��V��~u��i��V�^Wa?�����h�b�.��Vc�)H�Db]��05���ɓcp|�yU�_W.Ǆ�`��WD���WxDS�-�U�.V���%N���hɋ�P��� ʒ`lJ����ONr��Q����?����%�_&˿);VE�z�_���7�R�	t������H?�ř@$��K�7}ر9')�K��������+Z?��`I!�Jp���"�@pE��uz�L����j��.��ksu $!�Q��	����	ЀCKq���9��J�D��*����/��K�7��_��O�P������iֳ|SҦy��Ȉ�ݿ�9�"{����Cn"��q��\f�t����X��S��Dq��i��"I�JV�us��P��&�I�w���Z�tI�4���?v���҆Ef���Uґ�%�s'��.�qP�j�rsV;�-�wݱC�۹���}�Hr��MEf@vX�Oރ[|�7b��}nTd����U|�S�t�->*�[,��2G#(���k�T�UƘ�>����#�M7�犾����k��V��������rE�>1O���{H^�	>�gʧ^߻t�	�Wwz�h]z�Td�eYgAq��Q|U��%�Y�6[�� ��(m<;�fo�1�/s1d)�F=�|�<w�(D��"�k���*�����/PGO~��A�.�[���}�*�຃Y�1�Z�g�;�=�ל6�pe��"(;3�i��=���4/wy5����@��D�
�=��c�P@	�4V��'$,!�ע�U�.��ޫ|���KC�P]�P�Կx�����ר��}��w�b���ĹCF���UCn��Q�/���T֗N_�Y��,�qx�$�d�h��l�Ξ�=�.��]M3b�N��CP,JF������6Ւ
��p���	�$��^��Ƴ��NW���5�H�UCK���ǡ��Y?Lw�p_Lx���d �刀R[ "��)L���YgJsnO@��VI��$o_%�:X��J��rYm
^n����Tv�Ti�dc�I%���sȥJTH5Gڟd���x�c$�n�EJ�t�pȜ�/R����t��bk��Va�v־���y�2b�i�p�[���D9�o���m���
�ζ�Uy(��Ew�Mw�����[�5;��Vٛ�7ޙc���ߨ��8�
y�π\x`��]8&^&V���/_���xV�سT�ޙ�(FT�}���@h�2{����yD�/�	$	�rܥ�A+ͷU����x��|^<�����k2%�z�7=1T�r����,îӌ��J�^T=: ����yY��	�0�>*8�#�W`eٕ�}g��7���~�̦�3#����l��E׫u|�R�k]�?���}}&���R�*��ף)(��V�gpbi����wcu��+�[�4�r��Q{`U+Xc��QE����{U�{�t��)<�U^p���
.�F����(�6�j-���>��'�1�o�0�����e8H��=q�=��
}餀l�Z�t=7ƴ�O���w6�>�c�ʝ�eQ����:k�����b�dŚ��-�TB�UO ���x}�2yk2A�ȗ�8����*���;�Kvz�d��ypͳ�L7$����My��<�5c��m1^�4�6��������~� �1U5�B"^��H�����0A ��I�Ú�YF,�̹5!liw���������gl$b;�<��K^|L�}w��S�_�]����+��e�PEc_���ҳ9�:w�l��Rj���?��.{T�1(�e:'ٳ�e�:�Q���Y��p�x���[01E��
�G(U�j�����w�;<.Hʛ�����Xj�b�;a��Ao�R�����7�uz�ox7�����Q�����i�I�)�g��U��K!�p=�ps��M��8�;0Pp��"	�©DU����XT���r0���0��a�@=hΜ�����E����j BWN�~��C�w�T$��B������u?��!4��!O���V���t��(�ա�;RtE[?�3}ֹV�����HE�L�1� ��.�UqdN҉�.�aZ������"(���>�B�詾-���i�O�au�:���#8,!	!Z��P�Kx��~����xY��́XY ��Z`��ɥH�1������in.�A$��FO� 9���ܢ�����qS~n���!<���7����p� ެ�Lh�Q�w���Ӹ7�&�;��8~��[ѰvHd��N^�T��'�G�ɯ���RH�x�h�;�H )QYy8�B����j�n�8��m�$d3w��93�~�U���ۦݒ��F����PM���Kڗ��ɑ�ՇH��c
�	��d�gpLJ����NP��->/�سy1䀓����ٯ0����n}�!��曏�Ry�u�^|ir>�5��h���(ح�A; �T�y�/@�	_��0cr�w���+���|�R(|�	� �-ٮup��<���P�!X���&ѿkb,,�[�G�z)f���9jc�*��b�^&��ͿVDİ��9�W�Q���=���e3�)}C>��G��s�.~��	ˋ�E�O^�)����ӨW�6����<�VK��3��NDPc�F����S��f�������G5S� u&��y�����߳��P��1���7�*��)Q�3\�O�.��O���
�؍;�B���R��$C��vO��bb[����t��{��Z�7���*����,�w ;B���3�ze;E�b��X\ӧ&'��"���z���: �aJ]��2�kr����`����W6³@�p[*G���O�`�(�Ɵ�o��-'��m���D����r�t�]�\�H��b���r諝8��i��V:�s��;i$���L|�f?ffj(��_\��v���E���;�;� �H+�ABx�0N}𐥶�����N͇��r�Oz����F�!t�0��8�?c,:��c�`v5�,?���|�;ۛ��X��C�ӹ�B�����:�{����;o���8�����1k<*�VH
�YU[�|�#^D���H�JX����aaOLw�����Ǻ��~
���B+lG���5H?Z�@=Q�γȵ��c�_A�O���.�;ʬ���s?T����ea�>_y��fT��b���{�q�1������0��1���%����L،���_���݌������d�@�)�K_���0Z$��1�G0~2����Z [�!�N�c�|��a��N�8�7m���q�q�����D���&�Ѳ��%G�������%}8���ތx�木�K�i����"��B[x�ͨ�}jI�L�<�b��Cr����`$� `�N}ƫ�}p��鿋x7/�[��#�	MC��lw~���[Fu���c�Ysr���6G�0o����Ba:�4�߃�\G��p�� "F�����F��e�c[�)�r =^P֖g��~�P"&�_"�y��?��^ᾰLf���������G���1z&
|鱯���jU[��qi��I��h&u^�z�H%�҉���}��t9��vc�ʋ?[;��I����f���VkZ�VˤWP\aqi��� �J= �)�E۾��Q��fy����m�/�<��,�
��_旄+.|t�,ISZt�;�׆�kP��"WG��dL���%�x�TC��O��s�%MJ�
��h�sN��J�;t���f'�Z}�\�־m����Ñ�s·O��'����a��\=�<�^�×�R���,��L/��2$�_���?B��԰��sm��dm-8�Ld����꛹1�����^[���<���6��} �2���,�-�� ��p7��H���f�%n����������Ы��j���D�����|�W%�?pԗ�m]|�g�k���~jW��8f`\�\	���`m�'���\���:v�-8R���ۏB�\71����p�{��]�fX����,t�Z״N� ��K=6�V�Wsz�)#�\���zR��t��)�ͭt���E���Wf����4L��"�U&�%��z}mB�\�E����+�b܆ُZ����!j�zi�|3`'�x�xF,�i����
���W.Хr�u@�)���a�Nб��� >vv�>���<=�����.z��%	y�l�䦐K��3G_�ϰ8F�6
�����M�z�����!�`�_�F���,$��[�0}:h�#t�Q!��8��Py��'T-\E>v�s8~�'D�����X�V;��QV���I�^mOL}��g�V�%{�z/;�`�x��I
Z�S��T;mKz�(1�cALO��J痫�e93��ߺ9=���X�qҜ>������u&�>�x��:�9X,��l�mŉ��?[�4�{���&/�����$��Zw���L�1{�
��2��C(�u�W���9��7�H Aן�"�I�;��|]��}��OJD��}��%7V�����2�A������#aE۠��4�\P*�� �*y凪%Ze��A�_����eJ`���z�"+/�l�thb�" ���/��7�Z�-	���&L��� HQ�"29��S;c�Z�P�J�B��%p��1�E����y�A/��$C�/��a�w�����=�q�Vz�zg������Bv�9��ؘ�cP��L�YQi��v��� ������Q�~��5.1̢�*X�c����YP Qo!ATL,z"�p^�bg�	�	��s��O���fH�������GoB��2��H�Pt�-�u��X�A���:"�����݅���x�hb���;0�`����;�%�{4k3'���f��1ӫ����]dXb�f�7��#�.�Oӏ'2����|<d����y�9䜷�:�8Ȥ�_��wg��\;�z� r��m��~��1K�Y���)Z��p5*�ϯr�R�yO����~#�qC�DB��`�nxv�J��o�C��CL�߁�@O'�.',#EQ �2�%���3�D�� ˆ�y<���!���A)��f?)<V+0�5S7>�6��BV���u9;ՃmB�-EM��q��Y�VvĶ:4���3ȧ���27%�s�yA��k4i��(�p�T�����˧\}���Y��Mꔿ��� ��������G.F"6��o����q��j�vi��m\�	�)�A`��3��[~������c�H�a��8A��q��F�S�����;_7>T*�v	K��� ���sn�\�f��y'#2
銃A|Z�vIѹP��K�d���y�y�u���o'�%w^���9J�U�3.rz_��J��JQ�7D�=���36v[FAk�{(��7�Yԓ���`�淽w��eU���fb4�ʛ��g.92�=�u�>
�>>X������Qv��/wg���<����zu-X�܈�ðDLz�0]�d
���	nW;�
��u&�K��՝��2Rk�0�Ha�u��.��u_]~0�7��A�"x����!�.��mh��������j�'�΃~�Ęs���×�X�5	��\r��ܰ���u����5ɐ3V�jb:T�R)4��?�I�������t</�
m���AY��[hs�l����ju:���T++G��_�2�m�w�#����g�6"a�LgH��Y�B�`��e���ʋ+�3�!��jzY�l�p����g�0� %yY6T���Xo6�O��8&�z�c�A�%��Nm�8�y�O
6	�Qɇ7�3!�����/��u�o�a�5��"���--)5ړ���j��3�:�� �1��VUc:�qP=���< ����8؊&{F.���֥���'jg�����גj9v��:��t,R����J�#��[�s4��=zǾQ���,����ɼ�Q�D�Bh��^���9�?a��^�d�Kr��$�,���7�G�#�}�H"�����ԥ���| �5`ފ+�fB&�M�\H^b�L
���*��M'�(�B�R���с�u!��G�˻މ4��u[�oQ����4a�q*��0�E{���ic�S����P8C�p5��	+y�c��W�#1�v�B68oxkR�<�>��lў{�����cpU��cbS�y�75�Mٍ�-�%(g��"Z)Y�X���fp' �Ƞ��&P �p̓���� pp,4���?��X�]��32@Ô�9P����hx�wI��@�]�
���{$]��XF`�-���A���6�C��"�B,���g og�"��郂�w�Vh�G/�j�^tG%Y�7`֚~f���Nx�5$Z�����Y�W^��i��㗘ۨ���a<�*�d����T��a��Z�Q*m1W$������\ӦHV�1���w�J��;]���d���*�������!��H��⧖Uµ���YժD���1�t��?�%����ύ%��8?�l�p�Au��g)�NHZU��ʗ-k�&Q�yN�i������
k��*��}��S�ye�$f%몬fnI9kR2W̸��
v�U�x���o@�~4�]����]��B�ƙ����`6K"Ѻͷ�y:� ȏZ��{��o6����IҐ�"l���nh\g��j��!=B8/.����ݠ���~����-�3�+�Wt�m�\��:��]9��U"T6k�FV���6���� xn��/aT� q���i:������ڽ�<�+ԡSx�p�!y�L&-P~!QO��nU�[��8B�@��b\���l(�R��N�̀��<ܝ�����8�X��Os8�rK31V΃m��_����c��bdU<��&9G�D�pC�d|��K��KVQ4c�$�^�`G��h	���r����/ϗ!\���z~pn�1g"�����%Hr�6�J�tY�C�$g+��B%�<|�~g�@�a�ަ{�b/NX(�@�l��9o�,�� ��E�n����Wx�Ga-?�7���8���s5�C�G;���TcX�����`�������V��W��c�X ��ۗ}�����h��3J��k�`nxM�i�%>�i�� ɟk�:�)����H ,����#�Z�3 �ɷ�����_W��%nպ�;��:�:�ۛ��7�6�<F�HBH l R�
��P�n޻�>�����F�+�Z�Φ|���.�h�|Y�-Վ��%�w��c�!R�xCib�%�8��\��,�2>j\_[��I�{�[�H�-�[��V�mk)�@����� �Y�36f�l9�4�AJ�@e�{�I�p����ۑ6� (�z��c]wMef ��1ۖ]���ؿ�t�ƚ����R�8���R�k�<��uu7Ċx�i����,�S��_<c�������s=�7H��!g.��G�jk��@�X2�X�ȳ��R4h�s'��]-Sz���3���h-���@�"k8gZO�r�7⽗l��d�8l�����;�1Q�!��I�Ң|G���Q��X�g��v��Z�Uqd�i0�z�'�t��C	�䤰����%�pf�Lz��LV���kw�ش7Ĺ4q����6%:9��w3�	���J#��r� ��/N�k���pl	�FΏ��˧x�{cMs!���܇��da�.x]�*'o�m����!�-"�UsZ��-n�İQ n
&�6�����w.(&Uuؕ�%Y�ᐶ!�fS/���L�H&b7�;�җ
�l:-7|�S���@4"�h������7:i���?����I���~o΍������p85#�Ѣ��✛�����ǃBB�~����j+|�:����В��Y�֧�"de��wȳ���˸�4/�79���J_w2��@�nY6oYE�!	�G�,�{ �b�h[E�7���-��Gg��O�1RMaO�j����E�K�jL���*�$��>�?0�rxE� ����*�7H�I!�]O'w�������de�R%+-��Xē/�}h�-s�KFkP�ǅ���-Ďwx�4��
����g��ˤs�A"v1f����ک�]㨜��c&t�݋C�x%[=��%b�h	is `-����窱��M��!��$pCg`�K[�Ew9f�;@����W�h�_A�nz�U��i��=$"(F:ւ�tֵ;scQU�Ow�эrX��:��+���䉊�܋��jŘ��4��%j��EI/�Negp�?�����>K�V��Փ8��^L>6�t\�;r��ѽA�� o�����Kʒ�KwR�4>�.Kj\��s�`������r�ɩ]�NB̌)�O����_AX7�rO��v�4��~՘p�rK��=���um�-��A��/(��t��#��X6�"��A�*㉪��7s���@S��ãI4Fpܻ��qk:���1�/����HZ���1���_�2i~�ia�6�s��|D�75����/�6����� W�TvŮ[�uw��3�����0b��*���?`�T����ox	�X���pp\��۩�����(�QA�|˯˺/e��;�#o��P���)n��{�5������E�]��ʿ_�%�����ٿ� �?6E����0ik��m�MI�x�>�A+��=�,�ϒ�R!����ꀥb�):�w���#z�m��KC��0Oۍ�Qi8+b:9B^I�'��B�1$E?��'Z�Ր���lX ��c!E����8���L��=�d���pɹ�`y�6T�v�y�L�S�a�p�ʩ����T�E/LW
�%���v�o����;$'������w|��1JZMԴ|W4+4��#)�_aQ)�X�dB�?�Ƒ���;0:)�^h�#�P�U��c�*�J�݆r��ΟQ*R�>�zcԡ��j)*�~��W��1��Mp6��m��#�xL^���Њ�b�a������������4����iW-�U}񽕴�/��S'4�|�v;Y�ɋc�-{�i]G4�ᢛ�0fbٓ��h��=1�4h�|K�GT�����cd�gD��|#>2I@�Tذ�*�7;lp�y)��{�r3ܡ���W*�KYE�����엽q��X�؇uz{-�P�ʖ�f�X
�f�͂X	fO�m���\��b�\����[���-F�G��,Y����i�Jci��آ��t���_��؈��;[��Զ{��n��G�R%O�� P���2}��ml�a�2G8�������L�d/���h$ϟ��X�nf1I�Kmg�)���G_�ce)�]f�в/���w#���8p~/�;F�X�a3��ޗQ)���t��
�"��~e=���уVF7�����2ʱ1��KzJ �t�g�%�r� ��1�Tˏcj�B7�W�7��Y��7P4�ة2|��6g|��u�[��Ji�na��e_!{>���ΐ�N�\��ʄ_!�
�p�/3P_7�G���y;�^�i3a{��Y~H��XR���:�r�rH"�A����Oqٓ�hg�w�Lӻ���4SHV�������Mm�b�ѥ�┫����n���-��Z���1����'�!�%�0���E��]b���}gK��os���)�e���g�ب�U5&4��l�-��|�XQ&�|#�p���N�M�����oM��?O���� ��@�����j�+-;6+����U��Yut�<E�{�R��8���A��r���#��$u�sv&3u&�͔�T������ �A@'���v�u1ka�gpE���}:�S���ӵ��ס���"�usl�P�#J�Uː�jN��ߖ���&��m���!Wټ�#ka+�)J�s�ļ����Hԍ�C|B�N����욼?ER?�h��i79~� ��c�A�τA����T�Y��H4��!*\>�Ϭ@���ړ}�<�G����`L�i�S��]��
?�l�dp�v;E�T���۽��E|&��^�̝f�Kbi���ȅL�����]�=�;�����fru\�t�SQ���O8#��!�nR�����]��<�`K��d�����?8IK3Y���^О�Х�D��..�]�O|$��;�@�W1ݞ��x��|�����ܛ�m��^s�#�Qk؟���h�f ���"v��nPm����	�u�S>�X.$oH����sj����*���S���-���d�^8���"(�a�7�?�ѷ�nU2ld� �S�6J�\�`���ǽ��BT#�CU~��>]�K
0u{7aŗR�K����}���:3cb�c{M���㬒`z�Yk��#gW�#��m7���ٳ�o��ZӖ�Y�Y��[:����c3'q�Te��g�;tEb���"�"R������{��;�P����0b:J�D��;�s�rK#�cǼ"֑�ɩ��/�W�uqK��\�+�{��Xc�M�2���J�0�U
O�N���f\/����%�����j�%��ϔo)�玏C�Nc�l�-s�^�e�n."MA�u�ƹg`|�}����۪��l���I;���mB��O�g8b����
�]W|��39��$OⅡW��ξ��d�1e�x���qf5t��[l�\�2�G���$yx��@Q/�(�O���(�wLŌ����̹�
�e�h�z��5
�
����I�q�*{�C]�!ʉ�3ʤ!f�n0�n<��SjR�?���ߩ7�`$I�2Fɂ"6qiH�P��wPix\���6�[�{�I4����n�%�1[��!��U�-"݃�,�|=f�|܃SZ0%��Q�M�'�-%���G�qk�8��:�&�ls���2����^�*�d������p� "ʕ�aD����6	8P�|���*��B�9��Їޙ���A�p �� �4(ǖ~CT��+i����$�4����(�=�*=$%�Ha��+����P	�Cc�V��(�K<�.��	�Ϋ��:d¹��l��Z!��t@��m,���*y���u����@��\)���C���I��K��6p�yo��n2��-udl�b߫��;�>Q$,Y��g�2��P����Cr.�V�$%�7)o��^kq���&" ��qJJ�����8�'�)����LL���WF7��(��m�n��_����Z�H�4��#���!#sU@Y>�@�!\e>5o,o`e�-����4��ɎB���d�U|�_��2���qɩ@f�nd*_�g�9_TbH�9�_�[���X�6���91��-���CR ��t1,R+S���E��c�+A�Fc�����pi�$���4chT�=Q�0U�W���OwW=��Ygd������z@������D� ��^W��)�w�P���FP�	�X��uB.r���33�*B��?o	�b��=����D��_g٘8�6u<f*f�H�-�"�����W;x�������cV�$��'8�����a���������S������QG�I���/򪮈C��{]q������f�5�:�ع�'6@i��c�;Ú!{<�$���PH�2�x�G$W櫥�%�e��6�|��9�M���L�����k6a�����{��O�b��x�N����?R^�O���bɀ��@VU�;e��4�w��T�ա����P��*K�mB���Z^w�s���2�y�C{��9�|�G����iz�l2cՉj>������񹈆D��;�ZH~{�� �*?��\[|��^鄹nD3�9�?�c��}b���ؐi7�mV�[��4�K2�>�4�ɭ|��P�9��`��A]���5�C׍������ .A��yC?�4$.P��.�3��0����[�=��y0��iQ����Ajb�-�{�2{���:mI��G�%MmD�g�/���]QS����ISj��r�0Ͱ5F��q�%V���-��88���>��w�t�'�����Y��"��,�w an�yqL��A�#����N���-K�" �����rW�Y�DǛZ�^�_I �u�g�I�����3s�� �׭�}~�>�>=�`q�W��F�VM���]��s޴k�B�Oe\��/�l|ۆ�;�����o�u�7z�cCT2�b2�eky��mu������(�zeq�x9�aK�Æ7�l�ZJ�U���Si��S�x�>V8���ci�b�2�H�ɢ� �6Z��z��I�3���t�on�,CyD���(K�z*ʢ6��נ�mx��7|��G�-���RY-"3�z��?���T�����û�@��/�jϨF� nw���L4�
��R��Zn�{�P�Dz��3��7�M�������0�Y>��snC���^�֬񗴥�a��yٕK��­�ͤ#�{�7
�P�/���8���u�UY;�_�_� nu_W\5�����oK-�,�PCZD�H��������殽�#��G�e�x��ឪK��O}k]bBMmb|�|�߾,��B,���Qj5���T�W��鄇Z�Xԕ;8���M�����p��*G�B�y����=O�`J�Ņ�C��\����ʔ�Y��jlU�V��T{��b"��Ɗ^r����x"��������:Z�.c�^~P��	.p�9佶�ʅ;�9%nւ\P��e����w
]���G�{��R�.���sq�$Qx����3�.��6 Ǥ���*����̇gI��Jem�(��p���h��P�7-4�ސ��R��K�cf��m�čY���oW�kTO�$<r2a�Ⱥ�Q��l��Z��3�m�)�몢����v���Th�{?�)0�)��,��(���#Eq��Ӝ�J�Y;����凅¥����1��<������d�c�P`
�*Z
������a
��B`ҏ���ho�e��]3tb��ҧQ.�>��	����c/p�y)/V�*�Nu[\Qp��:��98�:���P�A���4Y���P�Fy��x��^�ƾHC�{�Q�V� |�+�^��4�����L�:s�m��!��?��-ǔ�����e,�RH��d�1����U�G�#�B�s\Z���k�Eb���]�a.%j��%�PI�>�&ժ��}w��mnP>Kuq�g�J��,B	������I����>6J�G�����㑉u�������W꽟~^��G`PP��lj�iaԆbz��4�ya+PިL���j�)���Ͽ�aέȟ[�{P���U���j���[΢������ftExU��'���W��d�~$���w��#r�OG�]C�Ny�q9�oa�b�+�xp����~ 5~�����ld�����9�x�:��{d"�$��x�$�(ph��ʂ[��A�%����>�t�����U���k�`#>���e,���J��]��N����ԅ�Eq����-{ͣ��N�ޟ:?b.s�]�̓�J��A��*��|���ȟ`Ɯ�n*?����EJs	��q+��`$,I[��̽�⛣'�C�MX-F`�{�C��Uߝ%]���{On<��+�CNcSy��٪>?����	�s��U�E�u��%�}%�~`�I+>s��
�\�4��C$%��o6�ɱ\�٠��b?Bq�2�G��	��/<�)�F�k��q A�Q�g��+�h�G�=.���~����bB��h�d��!�fa��;����$8��0�g�0r�y��'[�ه��o��@�4/�P|�����&���t]�>2�ӓӛҷP�صC��C���g����ʻbLD�((^z����\���E���v�!�QI�6`J�T1��܂�j�o�s�CZB��sLa͹��T�8���ƙ{EM�U���ʼ.�[G�V���k;�t�D�$8!�HR�>�.i��|'�2-Kx�BMRzk� ���so0˼B��a.���f���1j)|���(��B�ʋ��4�3�p�}�&�~�ωsQk�a�b��G���<�b����$��#��DCLV���x�x
��l�"C`�~�����%�{Y���(��j����gx���'�������	�Z��HSh|$�"B:HY�M�-Z�?3
������	]�@�kq)�6���ˑwA+8 ���8S|����6]y��iﱙ\D+	l`r�/p�ۺ�]@���EW˵�z��b�:Ù/�\����f|��+��b��t�m�B����G��x<���#ma�>i.
?�v��y�}j{�����%��"��p�N7P���<����%hd�X�+�8��������S�@�h��0�X���q>�lt�W�ϖ���M�Ysgݧ�
G)�q�\"�ᙩ�j�N�ثY�6�-�$Q0媀�k�X���GZY��2$^*JN��F�w��+#���If����Xæ㲈�o���Si��0l$�My��4-�]�h���^�������Үo�1�O	N�!1�~O�.�m]u�`��]�	,�<�{Rsla�Nt�2X0C^�%���, �>�$�)vk�Ӡ��i23Y �s���7@�q]^Krd3s�T��a���� Rzr�����\�(���ϑ�\�A�O~�%�L !�!]��
��(~	jD-䦚�w�Lw��b�u⬎��=/�:�zJ� (������|�/�9�O�Q���+��8&w����/�P�^��-��#��e�D�Ά5hi5*���d�����������8,�NJ���s�j��\�<6ӳ�>;���º�Ьǉ��bB�H����(�/�?tG����x��㞬_Swu�SըG?�Q�DS#uw�Hg	�4��+#V��N�~%��s�O�Z*;��+^f������yj�%�%i6��Vgb��qYdb���͂�Z����JS�Y���9S	�2�����	& �pj�O�ryP��p�gף�3�z+Q��B �<N���"Ee����-���]rd+`��ͱ�"u�GcjK�`�!�V���.�:�\)a15j���=;��"�F\�Q��(�F����u�?����E(k�� eS��j�[�5H�Z�;��Z~���[���߄�J��	����;��Џ����1���L� ~���aj��d�Yc�9X2��q���i|�&�ܵ��*W�
�4����d���rg�:�%s��A٪-�Ԧ�g>�df�0�M
XJg b�/�몙�ñ�Tj<���}3���10Q�L�l�6T9O �_&�/w��*�@������">r�B5.�qz��!;^�+Cl��=�@Nb}0أ����J/y:_���`L$%������^<.\
V���r�5��%�d��H�4$�jr.��Y߆�_=z
��娭к̐���"@�"aM����D�I`��BzbSF�5K��Zi�'�2^�{Z��&�����Ț�gb��kS���1���� �Z�Ls��@o� cw�:�z�.�*^��
����>�ƙ|�4p���b�����g� o��9E����Zּ��M}In�1VZQ��踲5�)H�"�sW(�6�R�w��*Z06�jѕّ������o������c[嶨�w�P��!t�a�J��O/,�l��F��LS��`��7֪jPZt�U���|$ 	}��i� (�u�do���7ה�c^��S��`�Ɇ.���rmdr0(��[�|I�k���������������C꜊�]QPVYb���?������ui�O��BH��x�Q3�Y?}��'����������8�w9�]Z۫L�O�M@ғ�ߣs��o��1�U:	nYi�D�;���7a�h]��l�b��ǀЊ@��A#a9?x�lg1���j���6��S ��E�S~=EP�V�`��L�U�_�S����tS)��@nn|�%�
�AN-Ǥ_��98��	5��":������V�!n�3h��^nI��_mɖ�>��_�����,Z�?�P�~P�<魅�6Y0�ta��qڽ���uT}�A�����ф�b��0]�/��K$6��d�T��� ieb�r�HQ�=؈��]b�����F��q�	��j]���D��O�1�����, ���{�l��c\���p��8�q�$p1Gom�0��j��g���^ v�ZQ�	Ӆ(L�N�-��Z���)��~��P�;�(��^ u,w�Z�X�(���4j����j�8 jz��3>4�K h���������f��Du�LMla	$A7{:�Q��^�̟s��Ǆff���q��U�$݁�Up���6�D����Q7vx��|{~���M�k�L�;���0:8!�0������m`4�a�4��4���EPr�9��Κp�5xHF	C�Zo�'?�ޖ��t4i��h{#�+�A�&��r������]��՞>��u|6.�����|���Qrڟ U�n���u �F���Ƌ���5e�ݣh���TPg�(�LS�fD�B��B;�jJ&�
�;�t��� t������	����I �i9g�ṱǸŸ�?n�[)�n��{EaW>@��N��G������,����q t�8�I��M���3�oU��`�"6uAs��$+x�$	�y����=AܢҢ״8U�8&
�Z�(�y�b��4�9��˜~��0︃�"(�*��fL��Ά<�!4ﷻ ��t�������P��.� ڶ�n˖;Vʻ;y�l.Jˁ�2�R��,�](I�%<�����>F�����x�v��Io�I)W��Z��3u~�x�٦��R�m��x��֯bذ��}�ͥk��ԣ��$��>v*D9z�ڨ8��������w��Xm�jdM;��DO 	>��n�Ct��-��E�O,L�/&��Fm8��b��W�� v�)_@j���J�����L�����|Up�;�4�^��gF�벙)�~�f�O0���5�_�'@?gU�[��t�eU�������߹�I�Q�����	l�2c���lݲI�nNA����e��Xڎ�V���"���S���F��bD����h���V�
 �
i�·�]aBtt$t��Զl�����:�j�#��'W`\�iڶ�AƜS������'L
]�=ed6TRު���8;����r�>�NɦL���w�,k���V�6�Ӭ�J�F�ѴPh�H�9w�+9�(Ǘ���4�8���z9�V|���Y)5E��D����Qf>���F�&%n��,�3W��f�����֨ �>�V� �;f��K嫩|g�	�Y�@e=M;��L l\ݦ��Ye���ȡz�����	���L*d�qKr<�N��*����Ѳ�o���qX��� �MA���9�$51�0�F�Y�P�+��'ߓܾ|�^���4�����&cǖ<ߊ�r.����|,���D���B\ �m��t�꿅p��J@�>k�QBX
BN�����A���ޢ�a^�a<) �� ��Z\*XW����x�͉</7'>f;e7y8�Y�4�Ɇ�N�S�o�6�� ��d�`{y�9�WRa'�y�r�����z$�\O�n����'���E��0j����J��U|)�"�.�p�K��� ����ґG��g8�k����gqu ��4�� �->r#���y����`�	s��E�c3ϸ�������BS�b������C��c���G-�CfT�*��ƾ�d��⁼��C����B�
����8�a�单�7���%.�Y5W�&]�����Ʌn_Tk�12�k�Z��H���Ll��˔,絭��|h�q�j.l���v�2�����j�F��g���f��cƣ�.���yٹ	���v9�B��9i�0P�b�#�����u�-�_`z��e��5VFB�� 
��-��7���� ċ���vY��ظ�/Ι<��šKt���S>H����T�_/lH�˟���6�H G�g���A"0�*�#W�'�ux�w���L ���#�HZw��|�~�r�#������8��&�/`��A˭�6�S�X�$KY[��pd~�d�"�H�oi���	������P1�U�fw��Lz?^��]�0�=��K*�O	<�8N�c=�鍎J���lZ��V�pT�X>�%H��L$ }?u(�$�z�e
&7�]�t3�l�p�}hZ�v�W����}9GI��1 14l;>9��|�S���5��BH-�\7+d� 2?��s�o`��x��Y�T������y�s\R����Z���;�)��D�A!eŤV<���Jd���\~.���g�ض�C�"]�`�) x۴E��,g���k��37�s;�P6����������|`M�y6���\�f�n�۫�s^��t��[�rLۼ�17m�n�>nX0�l��g_7�B�]�K��im�hhL��ՠ�x��K�k��d�m�����y RD�}e�ꆶ��ϑHגP\k{����8�>֡�՝uy��5�88�ƪ���B�ט�0k��U�@X�Htk�4�V��G���9L��'r�_{��XB{m�Ľ�9�UV`�r����|�-9��OI��;��:1A����!���0�}�ݏ(j.J1�Zq�wL�r��7�:J��s�}�9�2]�M��g�+[�f���~���n���vNevZ�$w�(��2^>HG�=5���?�4�!���KE�~?^~�R+�"���8z���P�����l�X��I���n�5��n�f�d�}-gJu��L���X�/�}*U͡%�H�e��F����Ki�l�Ij�C���)	�G�=D^��|8B��+�;�c^r���G�i���5����'H
!8�3=e���g�-�pl	��j�,�/j�饒*Sz�C �_-T�h� ~9{4->C�����~�l׈J螚N=�Lؼ�Lo��6�u��a���ƈ��I���í�-��Jz'e%�,�Ѯ�xP�����;;�a{�ب�Ƭ�s ?=So���g��13;p���*!��m����3��8P�䂦�����LmAm��a/�5gD��t�f����Ĭ�=!���ibi�弻w��`1���ݪ`��?�Osd��\��p�����8�ë��IF�{���y�z#��-j�떇�쓔�nZ�Fgi'�]������7lL+0�IH!��^�Y�.Yƿ4��P���U���`�^��X�RTA�?�G�GE�)F��p�w���%�8�!��wb�	�y︼:�ig��'������P����c
��1�x���^����SZKr�sB�	�Y���*��D{J�w�:(���/A=�$Ų#���_��xB��h���%<1U�1?��H�Y�+Î�-�P��޵��4*��N�C
nB�D�؅����3��5�j���չ9t�v����z��e�D�/W��-
Nj�˧l��I�uh�c͓���N�zBG�^��':T0`:�����1}DW�H�I5��5��I+}�\i9@�>���)�gK�"!�V`y���*rv�7���X�j�1��_n����.`(�Ia�>�D>C����N�`׋lQ�ە����}!�)��:*}(�hU韹�zHܞd�!IkJ�H�p�Ž�/�I� �3x[Z)�!'f��Ki?�n�)1q�2��m(5�3�Mh	8`����D�'ܱ%�����@M<��ᙯ�V$�̷n"H4�ӽ�r����A�j�)�4��c=�W�
[�n�#ϳ$v'����!ъ��4P�:P������G��/�1=����jE�7��oz �������V�}5e�Z�+�Ci��.V�G��x�2o�.��ѕG�,��?N[�6i�C�N	A�,�w;gބ1s|a�ŷ����)��ƆQ��%�c���L�Y�r�˴o���i������QU?:"�i\���Ls3��?��wbb��P���xa�~ג26�_��
$U��lM�P�y?�p�4��ҌQ�6u"�S��Kc26rK�-���V�����T�Q���������|��>L�B�����;�^�ܻ �-�C�Y�@m�����~M����LF����o8�C��#;��'��<�+�|��69E5̲�sن�i�^i����z�I?�#�{5{�����o�e�b̵d�c��(p��C~���8�[�Y���dS�d!��e �5�M�~�8�����)� �ܹB��{�loɆ����o"L"vt ���>�ו?�,6t��D���˓�IӖ�ei��sf��sk-^�9��VL�>	Y+�܆F"���էF��3a@-������u��R"R�w�H�$�ې���$�.s���)���U&��ftS��ay���AY���U�"�;z��������a�6ǯ�:�qΚ�+?x���M�r��0BĔ/-o~�,���T��`�~��<�e���7�I���s�g/8Q/��5��i��q����a�	[��g�,�/�IjpJ�Ɲ�]w�?g�+�fzdZ�ٿY���������h�D-K�#6� 7w���a�֘5�*қb�m"E�}��@��f@����c~�Q�b+�����Xbb"�^L:J�AL�E�N/�ի��y�t�ђ2ijy�v������-&r3{�����M��m��K����F�NDYL�MH�B�<;�o�D��	��J���T��O���4I�]��OM��O���2�9[�"��H�$�@��Ɨn��Ap �8����Yك�z���)y���Km}�^+-l|�]��1���(/l��g6�=.�� 典A�8:�,��^q��q* �*Z�o����bR�̍E�	��̞���, ֬�S��y<�JfƉ�0NyP�K��J�o�=_{vo��{Ѹ�h���N�J�b�`|��!���[ZM)�moP���{^QkPYuyċe�k�JMG�&�A[Ƒ��R�	�7M�k3L���on��ѫ[�@�#����{[����gt׳�Cc��/��TY�Gc��<5 wka[�~��t�T�K1�"E����J��=�i7��/ep���L ����n�u@&�f��+-�m�|� '|R���$��M֪� (�w\Mm/-�5^��~�!+���{�t�lh#@G�$ N��c��+�|�t��vt(֡=�)Gf.���/ɻ@@�`i*J����tй�ݖ `F��Hn���������'�R6�iu�ы̗�`��q���q�[N��1Ĭ>QQ��⽡������zV���
ڹ�qv�C��`4��<��Sa�G��˶n	�����k�Z*��~P=욽-?;���{<�U?��#�4|s�i��@��y��?s�x \}���F���ab���Xl7�����o��109� C��8n�I�-��G��������}�ق���%���*K��������������8`������s�ne�;�)�IM˫� �h�א��7�������^A-v�n^i���$_�"͟�F��L�z�hұ���8ۉ�v?� ":�I�����דuLy�d��+�a�]3�h;�}������?�چV� \W�U��aoUѻM�Y�1�ջFFR]���I=*d���C�b�j�t���'���jv���0�w�6h�(6�K~t����!ܕ�>/��.��R��h����l,{Z�=��n��OX��l�u�}�C�P�i�!S+E��3e	J�A���:��ϯ���S�:�Ƽ0ƹ��p�ٔ�6"N�T�H�K9���/�2����*IAg��?�0��@�[CL��N@��9��\'Gs�z�G�m��
͕x�ǣ�b�0�4L�t!v����v���D.��a�Մ�O�ҁ�Za\�,~��$���{�!'3K q�8���OF^�Ť�0�J'�J��|����v��r�l�T���E�����.n@��0ĳb��Ԗ�����$��{ƃ�(nش��~�[r-P5aT�3y��4�ư'���H7�>��;e����h���l��&��4D{a�_�kҒ�Ce�>��O.�H2A���U��GA.�*�G�9��: �*�Ǭ
x�Н�?��II� 7������}�J�>��4����� J�g��k�����4�E����)�1�}Jt�aN�>v�t'���������ۣ-9a��oǧ��fİ��h2���0$`tU?Hj�����0�;&`�����&�j�)��dV�7�ã�>�D�&���R�m�Y���Y��&��oSl�b���x���\d��;����
ӓ-,z6��vE�9����ï.骔eY\��d�Պ(�8"�?�3L � ��X�&Ӌ�
�!�I	����&�P�4���������y~���ډ8�L�6��N��v�<O�-�I~�9��h:�Nt�I�>k�m�sMb#Ǵ��b�yh�Tkl��`#���pB[p+𹹑��?(g*j����ϑl��Y/}n���^��t�`,�ۣ�+̷�K�3y��g��#���|�2�k03x��L�����o��m @m:�h��܏�ޏk~���!C�r��$�����id�:��"}���B���n�Fx0�.��I��`�0�}{�:Hs�D���bǩ@��N����6��|�4j����F'nOd��/�BB��6#e<�m�hܣ�U���d��r䏐�eNN5��Gm���
��j26 ��06��U��P<O���Fl.7&�&r�<���X?�A{AB��B2�j�5��4�ݍt��"k�i�Y�����蔢|Na���H�zs@Q�(�I!���8.���wcYsp!d�	{��a�b�X�����Y�wt�N���#�$�S���O���:W������xT�|���8�9���u�_&ݬɤI��ڝ�+��s�J�5Χ����dn+����cy��鎎��e@a�G-�cVy��ϸW/2=�X��0�����l�%ٸ��F��x@�r�2��3�%f���ASg�5+4n�j-Ŀ8�����DW�f��"�-@��>��F�!
�:����Y���C3����h�����+��Xhx�Wcj�s�5V�*��+�j��H�~��g�O]t��$����aȦP2G!`5G�K�`�Պa,|j«�5hc�'���������o�E���jCD�+��ɜ��~��OrI�Wd���!8*�I�(CA49+��|��&1�B����%��}K��)���Yo�cv7�s�(
@<Z_&7��t'���VRUq��A��JӋ�%�3�\��;�����y�дC�ָQw��w�v,�$�"�w�r�:!��%F�Lx�@�ܵ�k�%����B���֚F^ɀC��[�Z����_�����5H;34@���	��^P�)����&I���~�H$��%&O��Z*kX�o_�ƌ}��H)��B:hK��D���`6G�Q��~��i}��	�we�+ ~:�s�a|B����79����떤���	qL�b��2//�QBE���U�->�ػ=�D���a@X+ǵ֮E'Vv�v;���u(L(��7�D��O8��P�į(�evFl4�W�p��u�S���xt{�V�R���v��U�ڛ�0���ۂXP�n,�"2��O�ߡ%�����bP��쇥~b����6�[%;eR�c�˳6�)ֽ�漙�hn��(�t��烖��'���Q����>�%c�8#,�5��G`�'|�u+����kn��f�CBNm�π |7F����ɚ�3��f_^nD>�~@���]�a�E��x�+I����m`E�.`R^3�������7�s?L�y�S�8��������b�J	��f�U�����F��jDh�^�m;�~��,H��Ety�\	�qi�ۿ�"��X_P�pW��%�Ux9�Z����̑W,"I�A��@���|�n`�l�~��A�4�juؘ0��8d��~h��0�A+p�[�f�c���2�l��*6���q_qƾ6�؄��ޮ��L�j�)�����_������E����kh��� F�� �+�黦�px��O~'ć��e��a8w Vi��m�0�Q#;�����Z6��YH�AQaK<���z�uB&i��|�"J�o�e��S��~�#?��'�L[P��~HB^�=����)�s���7C/{��P3�t�O��k�Ϭ���Գ�}��A�i��1u���E����4�F:Y����0G���Ւ~�M�0hZ��G`�i��m�eM~9�@�E�t�ٺ���7���:��5�_��Ab�[������+� w<�.�SO�}h��+!�A�t��g�eJ����0��c���>M\�|�K~ͱ8>��d՝�}� _o�Ξ�ǌfT�'�����PP�$���� )6��;=�#����F��Z՟��P�;����'��z�*������<�.��'�\��,"˞n��C��_0e��>��0�_is��kŝp§J��T1�
�������q�`2���ښ��v�f�w��*G�$%N`G�u�ꞯ�k'�����B;-[	��N����ؑ@v�r�s��U=aE{)���N�鏗�g�����=����-�F�ͷg�k�(�hf��hO���F��,ů�]0�o� /�4^�Ů��^MF[uh�d��a;��{P�L&p7��]��*Hz*$�}��Vy��`�a��i��G�.��2Qڱ�Zإ�G���$؜��X D6���<l�h��c����p��+��Q�z���~���(�Qa�2"rx�N��_��e�4J|F�-��ą�!S�W�_ftc��kwV�x|r�����.]8	?�)��O�5�Lʽ�z�,s�1���e�5!)6u�	������Qn����4�NP��$��8���)��|�kc2)����9�QӴ̮p�!Tjb/	<LR+ �V2I�& ����ӂI��+�~RzH�A��
_E�-�����Ax��*7c���}|?�_��H�.Z�Lm���ٹ(ݼ��e��� K����J��)S(�u((�����w���ŭG�:ÿ��f����h�FU�e.�]`�7m�?�����;�zlA�l�(lr�>|Bl��Q��dA�6SU�F��9%m�� �t��`������h�&N�d�v��6��0��|�'=�����&�|���*��cmB����M���H}�g�9ͭ��8<(��|"RrV�S�U�;����; ��*#wg�,��J҅�����Ja�G��3�_P���|lf�/w6=���qĸ2.��"aG�=�>ւ7�œ\c�����<r~�~�����e��}�`�9n���(��<��9��(_�*�C�'޴}n�xw�b�bPj�z2˻�c��W%�E���@EZ�{噦Ë%cBvh{76�^T��1�7n-��~�­6{�[��G����VR~�/z^('�O�r��z �u��I�)�N-s�+�����Ͻ�v�����z�p��^���BV�n�No��{ΐ%���/5u�<�(��^���f���XRO�W��ـ06���+'� A=�P���Ũ�jz���~��o���3abZ+��e���7���&��E퉚�4�;�l��=���d�,S8g���t_��_/j�@�5y��m��ޔ�ɸ��������O�Q6��A����M���x��D�R�A�NE���e.�m	s��Yg�)����V��"/~4]�>��3�s5q��)��3��`�h3������({3��A��5��W"�'����7�-��ee�/*�j&��ԋJ�����J�}��v���Kr���T�[��,K�Y1��|��v׎��j��E�{S{�=��jj=��m�|�&�	�Ա6nIǈ%��áOE�.�������R9���u��ǯ|E�6!�0]��+#��t1l=���T�87>	�"��SH]�^���>�6�����P�Z��S�� �D������0ǎ����7���h")_F8��( �\A���ʜ���@�qt�2 i|�d������,|S�����)��p��uu6��i��c{�ϫ�e.K%Q�s��scF��Z�����/���u޹!�6~pb����
I�-��ѓu�ƪZ���Kb97�~�gAe�J��k͊��G ��h��&���,}w���O��0:���׶�@���Z_6$.1ϛ9���9������YWNX.�e^�����a�1/v�bx�$��^}��{���1�S� r�����&��̝C�%�Nd)R�gXip��0XS�Ue[�W
;^1�_B�<��/�2�_�2�m�k�D# �����XKh�ﶤ����<W�{8�5`c��qB
���S#��/e}�����W{��k�I�7��!q�^�a��Z��́�`"��%\SɆ�	��,�]κc���ܗ���o���N���u�!�&��&�{0���3����z�Dՙ�RD4Ә+�Гf�J3��Y����3xE�����=K+�wʯgD�������x�l_���|ޅ�"/����s���F�1��I�4�}��Z��r��|��JS�ӭ�YV)�(������wD =�����P
?���j�����c5B:�(�0��>�e�Ѧ��h��mU�z�p��i̿耀�Ȩc#}ʩ���N��ESe>�v3���)Ґ��@O�w���雞�Zq�~D�	L�V�+�klU7TgQvLMgĐ��Jɿ��P���?l���L��aR�3�.`����c�Y��Y�p�����cd���gI�~��	��@x�Ӥ�UP��H0��u%�4|���dDȹ��r���`X4m3����A���l�<ѝM��	���F+�婢1��V{vCuƎ��V����}��6q�p�m���zb_@� ��j��v</��ޣo^,�rEK=c��s�I1������'��y��[�.�Hi����=��K#}�PF������D��ar;��;�\���U7��U���2� _�[���kC�D��fa���l����-�7������v��U�_:הt��ϊ��>XGr�L��wy?t+(�	��=�������G����(��ݷ��:�YS�51�=˛�7D�b�� �IY���v	��>�~�R�B#��Y��p��l��LB��=�,��U�3Q�Z]6G^f@&��G�@s
A�,_;Z����KZ���h+cεډ�]����P�V�K�� LI��q~	�o*X��t�M��cX���sk��Q��Ak��"w���l��e0Z�:��;���ު&4ʱn(�r���\"��A6u��O�u� �.�O�E]$?*�04͛_�0�.C,.�s+�L1���Cs\�0��U܌#AC��� ��5��p*���aꤼ������#�9�lZK�J�\���Q*z�q<�EQ1d�d0���Ri����n��2(���/dh����pC���[�����	�v�ő%vWW�)�%��ڥ�ժ��P(.�F�1Q4�7��I3�x����?�G��¥�!�4*T`y魥s��mW���)�2n}��=�{5�i�U��)�7{r��g�������).�Cq'H����6s[Z{M��}li��9�e�p5�YR�8����B�����uh2R�vm���[��fU+G�q�c�>k1��[Y2�������u �3>u�^CI�E�cǝp�G`���4~�4����=�+�/fCn���Ԧ)��7C�(�p�I�m]�`�4�Jq�!���#`,�u���:�S�Pe�>�t�I^�����hsh+
�{�U�&}��G&��bz���kmAB�I�H�lq��nn��> NM�`��ܷGk�ִ<*WN�^q�׮4�^�U/��ާ?�����Ե��0��55��=�`���u�OL϶Z����҃���4C �.����4�U�:�3�E��d��4*�؆�Y�r�KO���4j�/����~��s�k?^�7q�ֺ&��Ҩu��@�M���X#u/���6\~�hT;�{b|.[�]��X������$�zy�K/�GQ�"N����HQ�a��R"��
C�'᧵���!8�l:�i0֏�%��(Fn\Gځ<�c����Ȕ��ŕ�@�.m����{�@�Jי3���%�����&b��l�$�S����uw�n'~B�9թ�� �o�ΆWF��X^�%"F���t~[��d���W��ʔ0����M���G��!3p��4���M����y�_r3s�܎�Y���6j5չ�71q�B�2�0�V!��ӡ԰��Ty1Թ����޲N&66z5�Z'I��f�f�.�H��Ț.�Q���*j�����f���ͣw���+
^���Rɧ u��)�\���t���>$h�.�d��g�MJ��K���U�c�E���W=��*¬�9����?Xz[�<���y����ͳS�9�פJ\�zFd��X�G)w�4g�4V'i��z��	S�:l�A7PKn:-s�wsn�ev�:���
a�w�EA�<bS�]�\�����Jk�ní:�-΍���q=��J��b2
�������>�+b�S�q5�9$ӕU�ï�g�~�">�#	WuO�� �rb_
���I�~LC�JM|�dmb�����4I�%z�#�eo5vT�ͨZ�`����Iv��X�F��T�3���s������Ke#^��ogN|����j��(��9�1|�Qy$���u[u������*������'pYP����A(s�R�I%��_�eziQ��B-f�@���rT�IL��WN����1��zV���hq�i�ŋ���O���{Be�*��@�1��M�Ur�I*�f]f��y҉"!�a�^I�<���p2���;C�S����a=��l�	��X��)�q0{��/Gi�2d>�˾��;R�o����e��?TO����ډ�����J� �U�=C��^��:��[.�Kr0Mn��߆&,\��C}�:OaYPP�]��Kv���\�{_Yl`��v|�ֈseVݤd�W��:��5�)�t������߬&~��V��>�W�5��8�a�ǟ�������2��&P2&Y�!�"ut�KV�\�Ni�$���储=��T\
�I*q �g��^[#�����\ �.iJN�z^����	٠��9�!2d�q�6��E�7(ƆnB*����e��L�cbri��1R�����'@K�+���I����i\��Wa��`����Y`�״�� ߰��v��Tn���\\�6��@7_���e� �8�a�5Fu���7�9.~�ݙEӽ�v�l䠬�L�/O*Z�l��[y�WRW;VZ��06�uF�c��!�<;���ڻ5�M[1���"oi��a9���w�M�T09N1�/|X�/�����e�^���8!צ����H�P[*�C)��S�=fz!����,�V�j�����\�=BܫY�������V"ܹ�G~�������?�$q O���3��E�%Dʑ碮���7+x{%�S��P��&��u������/�p�E�mųB��RD������-��Q7���7����0�&������_������y��2��7��1M�-r��f%�B�֌>E�,� >��g�؝a�7gx�ҷ�8�?�Q�Ժ�IS�4�:x���e,���D&�"�
HEG�����ګ�ơ5�?� Ėⳟʛ�M�U%��wS�D5��\�/��6Ɔ
���$~qi�'��*�&��3�~��v�c�E���;��w���|)��+vSX� 
��S�i)�����JsiJ�%umo���\�֥�3 p��Ni�O�3�zjR%�A{���WRֈ��Dm���̯�i����Q�hGgA�������So��;l�i�M̯��H��5(�M�����Q�9T���`�:����ԁX��U�\�����
@r)kJL}a�톎�S� |��ld����X�2
������]�r8��.�nA�Y��3��^�_K<Z�"ېH>kƋ��?6.<�+P�8�EA�.6�o�Q�ѫ�H[?�-��:�R�t�~�G)w��MҒ�^�c%l^dTC��d?ʉ\>:
č�y�`���U�0��k