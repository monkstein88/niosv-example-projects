��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$�������Vy�E�x�>�v���,���Qԧ���)s$�:��Y�m���Ru�.}ƀ��h?q��%W
�|���rk�>�m���yb[|T������>}������D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���y&+�W���^�D2i�>�|���B��,<��\ ��W�~��O�?��K��<$џ_�!�ʙ�E�T�0�61/�S�3#�=r��v�Ow��e�x8R��1۲��A`�ʃv�x+aC_>&���l��Y�D����@�ǟ��18�V� V٣�3����B>������Hd�.}�{�b�#<�w$Y$To+��]�aB{�b����t�°�����j���O�~�-V�?�3Ux@��\�I&��U���T�� z��_3�P��m��_ u�d{�[ֶ�vl_�c�U�k��74{�[��P��*E��D�㬩�#eZE��!�\�T���g4�ً ]rr����L�f�@�y�?Y`�MiG��	�G��W�L��ν�/���+
�F�	Ŭ�{R�� |�e3qŠ>���|Rф�Q�\-��Ɯ~�2���F*"���{E<� �֣�i�#Q*�wb��n
��_vA;�X�AMW�ע}�?TS,�u�[[?�aӰ�g��N��N4b��)��S�'3]3�4�n{g��!���ǽ�:�+_y�i�B�[ƶ��&���$_F�$vC �����}���f$YL���N�:��_z��>�(<�.�W�K�Kh a���,�6�K��Op2��1�Um�3��{����=e�u[�#��FZSWO$�.="�i� ��9��Z�����ETTZ��P���m5�b�Dy]�)y"c�r��b����ζ�N�:�wQ#�܊5��LN��<��+��D��r���3Zb��~'���ga�ۣ{V,������'��o�K�H(3���m��n��@�d��W�.A.PpI��73�v�2n�>�\��D&�=�S�1��z�Okk�y�	iƣ�jmY��f�=�E�)�T=�:�@rlO��-��$,)����C�e��:O�3��Ć5:��H�7�~7�9����KΚgX����	N�w��\a@�{��y�<�E����ɛf=���VI���M�+<HC�ɫ=��3�P������c}�52[��"������k�]���b�N6O��Ni���Q\U�cx�`�O���r�������閌�b���{�5�+k��/�W�5��ggk�Pn�1�tOI��c�!�bM�\�W$��y{��~)qa�+��� �~_�B������x�҅�@�WG5G�7�p�n0~cW����XX=����Z�Ly.�=���q��ב8��Piق�>�H/8�s��e JɣOz�}m������U��j ��)�e��\"x�"�=�"��(���so ��+�.�d�h�)�3�� A����'TN�� �V0Y�����=�1���,���'��֯���Z4ƨJ�S1�]Q0�l�lUsh�jU�w`���lNau�<��)zN�=�t�w�g�<S���Q6��:w��<,*D4d���*x�7�������>������[;Y|6V�l�5B�O�!{|���h[Z%��y1O(C���FR��T�2�pZg	$VbޙH�19�^�JeG "�xt	�4h1;����wG5�S��j����N+3rr��[>�d���"^c���E71��4ٲ��D�������NPU�+�F��s*]���t���2P>�duT�����s+�vt!d!���LTH^�J�AW��G�܂0��4�*M��J~��˅B���Fq~�"�P�RJ402�l�p��
��Lg~��P�G ��O�����2ܑXQK��m���K.��I��V3���!|a��_�j�6	0�
��rM���=o�0���wG����W:��'SF���D<F�(b"+G�v

O��pl�Y�t=s,����?F~Э�w��p�-���{��
�y?�_��3�2��C9G8*�����?B�]��v�b�A	�b���@c���7	T����I�𭮋\p[��R/����p��d���J� t1��=����R�_��G����RCO��ۻE't�͠a?�W���y
l��������{7��~m`t[���3rFJI[�*{���Y���o��̋	l��|��L��j<��߇�*��w�W�u�P�Cܑwu���4\��hF.�~'����_����$x}*���&/�� ^~ ��g��k��o>�"�d�1V񏡴����T������H��O|���-����iM�eki�j��ݬ�yt3��v�k�X���K�j,a����t��B5���jZ����ef�փ���T�ߵ/�1�:�U�h��6��h��v.�\�Py
�ß��T���E��s����u2I��\73�.^\nJܠ$������?f[��t͎�EU�yʪ���~�_E\q�)�R
)��i����I����˵�Y��I��<�;̫������O���#����/��Y�d�/o���RuS�)�L�e�8��y<�Vğ�����C�]�/\�.��k���� �\�#���v=B�ܲ�lI�N��[�Q�?&���,�����,O�!b�A��҉�t����;��Cgǡ��^	�q�C�^�{�����1Y�����!;�).)@k���UV�:F7�J��{�g� �"���
彴G��ԕD�*%CSv��6"��t����$��1g���h L|
�5���Tr��l�Lr�d��a�(��E�M���#�%�RfZ�p�4���)i�	��=���&6�k�6����� 	z����]�SqLw ���ߵ�Eq�8�a�PI�~w�Bz��X�K�Uts�4����7m�͝s5��5��G����~�(�����V�M�vq���{V�3U��^��(3�/��Z��Mc`.�LAAY�qɔ��V�h���5���V.��ּyP����h�\2l�¿��8y<m[97��z`�;�?�pɤ�!��5��N��&��B�0�k�o/�Hz��	|�	���J@���W�ǻR�ۅwM�X�$zc��o�l���:j����	T�|٩¼ru��c*=v�-hX S�fMR�1io����J�y�sR�������hWhͣJQ��|����>����F�$����U�/I)�緓譈���K'�6�DR��3|��w���۱���.�J�|�fa*nS�$??6M�"6x��K��zo�*k�M"��ψI�����'�:��(�eQÉ!F.�H!�eܒp����Yv��_��.����&r����d}�aṦ�02�������z���XS�Uj���(�%s�1A�Y�ZT�})o,u		�����0��[�u��=�$A�����l���F�Ʃ�-���3{w�枌Sb��h��V/�8!�0��2/�-�^V�qـ;"""��={����H6���I�=�q���p�17sa���#F&�$j�6�V1,Ui�lh�HDde�y�eͯ��F��7b�g}��
U.���1�����!:&W��"$pn.3�ڙT,*��q��I�b ��H�����# �ǥ �"��(�%��}BY���Mܗ����&PB�����M�g�HU�@�������f�q�����k&��7� ��$j��~�>2a^���c��pep#�v���kTN��;���[��i�I��olR4ļ[ٰ� PT����&�On{�_��p(�l(�&'��1�cDe�����i����<a���㽦Nюr�v5�Q�F��u���Р���$�4ӣL��l�ϟ�<.]��/��N%���'��k���o੦^;:cZ�_�ʌ��oa}�f;�k���C��E��؇���;X���!)���k�ɖ�+�J\���T5��aخh�`FA�DV�V%y�6Ǯ��3��&����ă�Mjoݟ2�E�����%uN{�Ҹz��U�lt����q����7����@(&V��_�:R�Sۦc+��BH���%�@���v���D$Ŵ�҂�C~o?�� �v7L˴L��������;������j$�m,�sE#g�����4�?l�'�g��ߴ����z�C�r��j�'�]=v~�:��}{�I�^��2��emɱ��������f�%��6j6�AE��4YEj��w��l�vO����P;菺49EU���ط�V�5^�ڣn�ްm�f��
$3(��h�r�ׁ8���k�o�Z��w����
���9�cZ;�:����bԣ�W&i_�ElG�Y�Kw�~�ӹ.h�:�4K�w�Nu���=�&�,`��d����̧�|ƈ��g���A������G�d`�t�ڣC���>(Հ�ѩ�x�N�em��9dS��vJG���X}��c��7[mf�j��Ē�xBT��q��$3�
����7��j�a��֢˿2;���|O�����2*��g��ylbA��e$|��yx����Al*M|ֽx�7E͓����<l�9�_O����}Hg�q2��>�R�[�%��xo��i!G�����c�%�"6��.�N'ݍ0�����K����{P4�$�M�=6�8w���=�B�:m�C7Ӝ[>�L��w#<lQ����K�c��n���7�	�E�63-��&g ^�"keK����ָʡ��j�g�&Q�߱˚!����$��J�V+}�,��;�Cm& ����.�οL_xv�.�3���d&��	4�#C����dW���F��x�!j���]Ss�o/Ьl���;>����@�:&Zt�:$�Ĕ�Q�_>p��N0�@_htc��W�ReP8��7�<�+=Uo-��q�gz�72��ARX)���i�}@��q}~8��������]�|O��X��:!�裧i�ǆ|d��r�u[��췋[96�����@���D@q��1X!q�g�Xl@Fs�O��g1+R�TE&"1gܰ�������VG+g�b�? 9�s���A����pbNC�f#�N����6������F�s�&�C�n �ʞt��f%�{Z��f+��8Iشu؆%G�wZh��Mȉ��ċ�Y�&�*��t��[k�٫���m��>��t�D+ϑ>���h8����`��S�pS�	�f0G�;@w>��Oۭm69�};���I��ah�'��&�@��j�tQ�=w$~%e;W[>{z�� S��;���L����@ ��$b!:u��6���]9��du����߶���D���ś�ϼ�;5��L�jo,�:{$\��E.��B��\f:ܪg�z��5c�����	���GB�� �� p&Ɖ�񖬒�R���i��K�?�P\B�������{` �Z�����AzxOdr��cay)>@7�/�mVU�J-��������7��T��3�K �:8�I���SW`p�j���j&՛)x-a������pǞ���c���h�vwe�Xе��~�Aٜ��30�j��B�����v Ӝ��ѧ>�"u#�U̲%	���E�_�f�b �:S�^��[>�g���kP�b8�7�<bV`��'���Q�U-�������$1�!��oP���v��bD�OW������2y0��O��B��x|<�O�s�ۊ:�H0T���/�����.�%���3�^�{{�78�}���p��_
O�K���t^@><KVWC�C�:�����W*?N��dK�TI6�:K%������k@=��9:(���p��21��翤_�1�MJ�?	U���mr��FJg�?��\eX�tذ����s��T&h����ڟ��5��9,�L%r��I��TF��Hzu�ߛԿ؝� 񩺰f��#�,4�
��#ִ�����,�i��5��9�5G������>�����^ ���t����6��X��'�ʯ3HJ9�^V�k���Z�<�h�����;�Ų��G &������g������������a�����a�hu����@S��H��q���._9T���ͪ�*i)C�Kdn�bkA��C�M�u�ϳ{�	��P]��C�2�dC�#D���+J���7�J[j�z���wj:=4�/��������g��f�ToP?��Z�r������ulay/$�?D�ף�+eMp���]�� ���$�"�SVr;.F�>:���9�F:��*�~3_l̶,�X����a��yT�O3�H�<��^9C�z�e1�=%>e�# � *G	-�_!T#��B1b�b �NB��A�&̭fd����`P��Xi��#<F�5ۍ��k��e�{�~=��9Φ)6��/�b��b�O %�0$�[�|s�r�Hs|Ѫ�kO���I%Q&슠�D�J��ɨH��	���g:R6��aypV�ނ���,��z'�r���B]�?ݲ��z�ځ��e���Y�1an촯�I�&�w��)�=\݋r�	v؅U,+~�8�5�c:�b72�q;�E �2�n��ʉ���%VAON�k3G}	�u"�X�`�N]`�ke��~U5u���8o��Cwf� �Y��v���f�{|8/x����vgV���aɤ����Q��qƨ�����?Ѓ���\~-���b�8�jg�u�h��?�{��jK)�$�wd.����`�q�P�����.�zTO	��0�E��).��|�k6wMBd���㯼w�!%�R'���==�����r8�����S:���Z�I[��O